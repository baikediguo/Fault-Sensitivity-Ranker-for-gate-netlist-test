`timescale 1ns / 1ps

module tb;

  reg \A[0] ;
  reg \A[1] ;
  reg \A[10] ;
  reg \A[100] ;
  reg \A[1000] ;
  reg \A[101] ;
  reg \A[102] ;
  reg \A[103] ;
  reg \A[104] ;
  reg \A[105] ;
  reg \A[106] ;
  reg \A[107] ;
  reg \A[108] ;
  reg \A[109] ;
  reg \A[11] ;
  reg \A[110] ;
  reg \A[111] ;
  reg \A[112] ;
  reg \A[113] ;
  reg \A[114] ;
  reg \A[115] ;
  reg \A[116] ;
  reg \A[117] ;
  reg \A[118] ;
  reg \A[119] ;
  reg \A[12] ;
  reg \A[120] ;
  reg \A[121] ;
  reg \A[122] ;
  reg \A[123] ;
  reg \A[124] ;
  reg \A[125] ;
  reg \A[126] ;
  reg \A[127] ;
  reg \A[128] ;
  reg \A[129] ;
  reg \A[13] ;
  reg \A[130] ;
  reg \A[131] ;
  reg \A[132] ;
  reg \A[133] ;
  reg \A[134] ;
  reg \A[135] ;
  reg \A[136] ;
  reg \A[137] ;
  reg \A[138] ;
  reg \A[139] ;
  reg \A[14] ;
  reg \A[140] ;
  reg \A[141] ;
  reg \A[142] ;
  reg \A[143] ;
  reg \A[144] ;
  reg \A[145] ;
  reg \A[146] ;
  reg \A[147] ;
  reg \A[148] ;
  reg \A[149] ;
  reg \A[15] ;
  reg \A[150] ;
  reg \A[151] ;
  reg \A[152] ;
  reg \A[153] ;
  reg \A[154] ;
  reg \A[155] ;
  reg \A[156] ;
  reg \A[157] ;
  reg \A[158] ;
  reg \A[159] ;
  reg \A[16] ;
  reg \A[160] ;
  reg \A[161] ;
  reg \A[162] ;
  reg \A[163] ;
  reg \A[164] ;
  reg \A[165] ;
  reg \A[166] ;
  reg \A[167] ;
  reg \A[168] ;
  reg \A[169] ;
  reg \A[17] ;
  reg \A[170] ;
  reg \A[171] ;
  reg \A[172] ;
  reg \A[173] ;
  reg \A[174] ;
  reg \A[175] ;
  reg \A[176] ;
  reg \A[177] ;
  reg \A[178] ;
  reg \A[179] ;
  reg \A[18] ;
  reg \A[180] ;
  reg \A[181] ;
  reg \A[182] ;
  reg \A[183] ;
  reg \A[184] ;
  reg \A[185] ;
  reg \A[186] ;
  reg \A[187] ;
  reg \A[188] ;
  reg \A[189] ;
  reg \A[19] ;
  reg \A[190] ;
  reg \A[191] ;
  reg \A[192] ;
  reg \A[193] ;
  reg \A[194] ;
  reg \A[195] ;
  reg \A[196] ;
  reg \A[197] ;
  reg \A[198] ;
  reg \A[199] ;
  reg \A[2] ;
  reg \A[20] ;
  reg \A[200] ;
  reg \A[201] ;
  reg \A[202] ;
  reg \A[203] ;
  reg \A[204] ;
  reg \A[205] ;
  reg \A[206] ;
  reg \A[207] ;
  reg \A[208] ;
  reg \A[209] ;
  reg \A[21] ;
  reg \A[210] ;
  reg \A[211] ;
  reg \A[212] ;
  reg \A[213] ;
  reg \A[214] ;
  reg \A[215] ;
  reg \A[216] ;
  reg \A[217] ;
  reg \A[218] ;
  reg \A[219] ;
  reg \A[22] ;
  reg \A[220] ;
  reg \A[221] ;
  reg \A[222] ;
  reg \A[223] ;
  reg \A[224] ;
  reg \A[225] ;
  reg \A[226] ;
  reg \A[227] ;
  reg \A[228] ;
  reg \A[229] ;
  reg \A[23] ;
  reg \A[230] ;
  reg \A[231] ;
  reg \A[232] ;
  reg \A[233] ;
  reg \A[234] ;
  reg \A[235] ;
  reg \A[236] ;
  reg \A[237] ;
  reg \A[238] ;
  reg \A[239] ;
  reg \A[24] ;
  reg \A[240] ;
  reg \A[241] ;
  reg \A[242] ;
  reg \A[243] ;
  reg \A[244] ;
  reg \A[245] ;
  reg \A[246] ;
  reg \A[247] ;
  reg \A[248] ;
  reg \A[249] ;
  reg \A[25] ;
  reg \A[250] ;
  reg \A[251] ;
  reg \A[252] ;
  reg \A[253] ;
  reg \A[254] ;
  reg \A[255] ;
  reg \A[256] ;
  reg \A[257] ;
  reg \A[258] ;
  reg \A[259] ;
  reg \A[26] ;
  reg \A[260] ;
  reg \A[261] ;
  reg \A[262] ;
  reg \A[263] ;
  reg \A[264] ;
  reg \A[265] ;
  reg \A[266] ;
  reg \A[267] ;
  reg \A[268] ;
  reg \A[269] ;
  reg \A[27] ;
  reg \A[270] ;
  reg \A[271] ;
  reg \A[272] ;
  reg \A[273] ;
  reg \A[274] ;
  reg \A[275] ;
  reg \A[276] ;
  reg \A[277] ;
  reg \A[278] ;
  reg \A[279] ;
  reg \A[28] ;
  reg \A[280] ;
  reg \A[281] ;
  reg \A[282] ;
  reg \A[283] ;
  reg \A[284] ;
  reg \A[285] ;
  reg \A[286] ;
  reg \A[287] ;
  reg \A[288] ;
  reg \A[289] ;
  reg \A[29] ;
  reg \A[290] ;
  reg \A[291] ;
  reg \A[292] ;
  reg \A[293] ;
  reg \A[294] ;
  reg \A[295] ;
  reg \A[296] ;
  reg \A[297] ;
  reg \A[298] ;
  reg \A[299] ;
  reg \A[3] ;
  reg \A[30] ;
  reg \A[300] ;
  reg \A[301] ;
  reg \A[302] ;
  reg \A[303] ;
  reg \A[304] ;
  reg \A[305] ;
  reg \A[306] ;
  reg \A[307] ;
  reg \A[308] ;
  reg \A[309] ;
  reg \A[31] ;
  reg \A[310] ;
  reg \A[311] ;
  reg \A[312] ;
  reg \A[313] ;
  reg \A[314] ;
  reg \A[315] ;
  reg \A[316] ;
  reg \A[317] ;
  reg \A[318] ;
  reg \A[319] ;
  reg \A[32] ;
  reg \A[320] ;
  reg \A[321] ;
  reg \A[322] ;
  reg \A[323] ;
  reg \A[324] ;
  reg \A[325] ;
  reg \A[326] ;
  reg \A[327] ;
  reg \A[328] ;
  reg \A[329] ;
  reg \A[33] ;
  reg \A[330] ;
  reg \A[331] ;
  reg \A[332] ;
  reg \A[333] ;
  reg \A[334] ;
  reg \A[335] ;
  reg \A[336] ;
  reg \A[337] ;
  reg \A[338] ;
  reg \A[339] ;
  reg \A[34] ;
  reg \A[340] ;
  reg \A[341] ;
  reg \A[342] ;
  reg \A[343] ;
  reg \A[344] ;
  reg \A[345] ;
  reg \A[346] ;
  reg \A[347] ;
  reg \A[348] ;
  reg \A[349] ;
  reg \A[35] ;
  reg \A[350] ;
  reg \A[351] ;
  reg \A[352] ;
  reg \A[353] ;
  reg \A[354] ;
  reg \A[355] ;
  reg \A[356] ;
  reg \A[357] ;
  reg \A[358] ;
  reg \A[359] ;
  reg \A[36] ;
  reg \A[360] ;
  reg \A[361] ;
  reg \A[362] ;
  reg \A[363] ;
  reg \A[364] ;
  reg \A[365] ;
  reg \A[366] ;
  reg \A[367] ;
  reg \A[368] ;
  reg \A[369] ;
  reg \A[37] ;
  reg \A[370] ;
  reg \A[371] ;
  reg \A[372] ;
  reg \A[373] ;
  reg \A[374] ;
  reg \A[375] ;
  reg \A[376] ;
  reg \A[377] ;
  reg \A[378] ;
  reg \A[379] ;
  reg \A[38] ;
  reg \A[380] ;
  reg \A[381] ;
  reg \A[382] ;
  reg \A[383] ;
  reg \A[384] ;
  reg \A[385] ;
  reg \A[386] ;
  reg \A[387] ;
  reg \A[388] ;
  reg \A[389] ;
  reg \A[39] ;
  reg \A[390] ;
  reg \A[391] ;
  reg \A[392] ;
  reg \A[393] ;
  reg \A[394] ;
  reg \A[395] ;
  reg \A[396] ;
  reg \A[397] ;
  reg \A[398] ;
  reg \A[399] ;
  reg \A[4] ;
  reg \A[40] ;
  reg \A[400] ;
  reg \A[401] ;
  reg \A[402] ;
  reg \A[403] ;
  reg \A[404] ;
  reg \A[405] ;
  reg \A[406] ;
  reg \A[407] ;
  reg \A[408] ;
  reg \A[409] ;
  reg \A[41] ;
  reg \A[410] ;
  reg \A[411] ;
  reg \A[412] ;
  reg \A[413] ;
  reg \A[414] ;
  reg \A[415] ;
  reg \A[416] ;
  reg \A[417] ;
  reg \A[418] ;
  reg \A[419] ;
  reg \A[42] ;
  reg \A[420] ;
  reg \A[421] ;
  reg \A[422] ;
  reg \A[423] ;
  reg \A[424] ;
  reg \A[425] ;
  reg \A[426] ;
  reg \A[427] ;
  reg \A[428] ;
  reg \A[429] ;
  reg \A[43] ;
  reg \A[430] ;
  reg \A[431] ;
  reg \A[432] ;
  reg \A[433] ;
  reg \A[434] ;
  reg \A[435] ;
  reg \A[436] ;
  reg \A[437] ;
  reg \A[438] ;
  reg \A[439] ;
  reg \A[44] ;
  reg \A[440] ;
  reg \A[441] ;
  reg \A[442] ;
  reg \A[443] ;
  reg \A[444] ;
  reg \A[445] ;
  reg \A[446] ;
  reg \A[447] ;
  reg \A[448] ;
  reg \A[449] ;
  reg \A[45] ;
  reg \A[450] ;
  reg \A[451] ;
  reg \A[452] ;
  reg \A[453] ;
  reg \A[454] ;
  reg \A[455] ;
  reg \A[456] ;
  reg \A[457] ;
  reg \A[458] ;
  reg \A[459] ;
  reg \A[46] ;
  reg \A[460] ;
  reg \A[461] ;
  reg \A[462] ;
  reg \A[463] ;
  reg \A[464] ;
  reg \A[465] ;
  reg \A[466] ;
  reg \A[467] ;
  reg \A[468] ;
  reg \A[469] ;
  reg \A[47] ;
  reg \A[470] ;
  reg \A[471] ;
  reg \A[472] ;
  reg \A[473] ;
  reg \A[474] ;
  reg \A[475] ;
  reg \A[476] ;
  reg \A[477] ;
  reg \A[478] ;
  reg \A[479] ;
  reg \A[48] ;
  reg \A[480] ;
  reg \A[481] ;
  reg \A[482] ;
  reg \A[483] ;
  reg \A[484] ;
  reg \A[485] ;
  reg \A[486] ;
  reg \A[487] ;
  reg \A[488] ;
  reg \A[489] ;
  reg \A[49] ;
  reg \A[490] ;
  reg \A[491] ;
  reg \A[492] ;
  reg \A[493] ;
  reg \A[494] ;
  reg \A[495] ;
  reg \A[496] ;
  reg \A[497] ;
  reg \A[498] ;
  reg \A[499] ;
  reg \A[5] ;
  reg \A[50] ;
  reg \A[500] ;
  reg \A[501] ;
  reg \A[502] ;
  reg \A[503] ;
  reg \A[504] ;
  reg \A[505] ;
  reg \A[506] ;
  reg \A[507] ;
  reg \A[508] ;
  reg \A[509] ;
  reg \A[51] ;
  reg \A[510] ;
  reg \A[511] ;
  reg \A[512] ;
  reg \A[513] ;
  reg \A[514] ;
  reg \A[515] ;
  reg \A[516] ;
  reg \A[517] ;
  reg \A[518] ;
  reg \A[519] ;
  reg \A[52] ;
  reg \A[520] ;
  reg \A[521] ;
  reg \A[522] ;
  reg \A[523] ;
  reg \A[524] ;
  reg \A[525] ;
  reg \A[526] ;
  reg \A[527] ;
  reg \A[528] ;
  reg \A[529] ;
  reg \A[53] ;
  reg \A[530] ;
  reg \A[531] ;
  reg \A[532] ;
  reg \A[533] ;
  reg \A[534] ;
  reg \A[535] ;
  reg \A[536] ;
  reg \A[537] ;
  reg \A[538] ;
  reg \A[539] ;
  reg \A[54] ;
  reg \A[540] ;
  reg \A[541] ;
  reg \A[542] ;
  reg \A[543] ;
  reg \A[544] ;
  reg \A[545] ;
  reg \A[546] ;
  reg \A[547] ;
  reg \A[548] ;
  reg \A[549] ;
  reg \A[55] ;
  reg \A[550] ;
  reg \A[551] ;
  reg \A[552] ;
  reg \A[553] ;
  reg \A[554] ;
  reg \A[555] ;
  reg \A[556] ;
  reg \A[557] ;
  reg \A[558] ;
  reg \A[559] ;
  reg \A[56] ;
  reg \A[560] ;
  reg \A[561] ;
  reg \A[562] ;
  reg \A[563] ;
  reg \A[564] ;
  reg \A[565] ;
  reg \A[566] ;
  reg \A[567] ;
  reg \A[568] ;
  reg \A[569] ;
  reg \A[57] ;
  reg \A[570] ;
  reg \A[571] ;
  reg \A[572] ;
  reg \A[573] ;
  reg \A[574] ;
  reg \A[575] ;
  reg \A[576] ;
  reg \A[577] ;
  reg \A[578] ;
  reg \A[579] ;
  reg \A[58] ;
  reg \A[580] ;
  reg \A[581] ;
  reg \A[582] ;
  reg \A[583] ;
  reg \A[584] ;
  reg \A[585] ;
  reg \A[586] ;
  reg \A[587] ;
  reg \A[588] ;
  reg \A[589] ;
  reg \A[59] ;
  reg \A[590] ;
  reg \A[591] ;
  reg \A[592] ;
  reg \A[593] ;
  reg \A[594] ;
  reg \A[595] ;
  reg \A[596] ;
  reg \A[597] ;
  reg \A[598] ;
  reg \A[599] ;
  reg \A[6] ;
  reg \A[60] ;
  reg \A[600] ;
  reg \A[601] ;
  reg \A[602] ;
  reg \A[603] ;
  reg \A[604] ;
  reg \A[605] ;
  reg \A[606] ;
  reg \A[607] ;
  reg \A[608] ;
  reg \A[609] ;
  reg \A[61] ;
  reg \A[610] ;
  reg \A[611] ;
  reg \A[612] ;
  reg \A[613] ;
  reg \A[614] ;
  reg \A[615] ;
  reg \A[616] ;
  reg \A[617] ;
  reg \A[618] ;
  reg \A[619] ;
  reg \A[62] ;
  reg \A[620] ;
  reg \A[621] ;
  reg \A[622] ;
  reg \A[623] ;
  reg \A[624] ;
  reg \A[625] ;
  reg \A[626] ;
  reg \A[627] ;
  reg \A[628] ;
  reg \A[629] ;
  reg \A[63] ;
  reg \A[630] ;
  reg \A[631] ;
  reg \A[632] ;
  reg \A[633] ;
  reg \A[634] ;
  reg \A[635] ;
  reg \A[636] ;
  reg \A[637] ;
  reg \A[638] ;
  reg \A[639] ;
  reg \A[64] ;
  reg \A[640] ;
  reg \A[641] ;
  reg \A[642] ;
  reg \A[643] ;
  reg \A[644] ;
  reg \A[645] ;
  reg \A[646] ;
  reg \A[647] ;
  reg \A[648] ;
  reg \A[649] ;
  reg \A[65] ;
  reg \A[650] ;
  reg \A[651] ;
  reg \A[652] ;
  reg \A[653] ;
  reg \A[654] ;
  reg \A[655] ;
  reg \A[656] ;
  reg \A[657] ;
  reg \A[658] ;
  reg \A[659] ;
  reg \A[66] ;
  reg \A[660] ;
  reg \A[661] ;
  reg \A[662] ;
  reg \A[663] ;
  reg \A[664] ;
  reg \A[665] ;
  reg \A[666] ;
  reg \A[667] ;
  reg \A[668] ;
  reg \A[669] ;
  reg \A[67] ;
  reg \A[670] ;
  reg \A[671] ;
  reg \A[672] ;
  reg \A[673] ;
  reg \A[674] ;
  reg \A[675] ;
  reg \A[676] ;
  reg \A[677] ;
  reg \A[678] ;
  reg \A[679] ;
  reg \A[68] ;
  reg \A[680] ;
  reg \A[681] ;
  reg \A[682] ;
  reg \A[683] ;
  reg \A[684] ;
  reg \A[685] ;
  reg \A[686] ;
  reg \A[687] ;
  reg \A[688] ;
  reg \A[689] ;
  reg \A[69] ;
  reg \A[690] ;
  reg \A[691] ;
  reg \A[692] ;
  reg \A[693] ;
  reg \A[694] ;
  reg \A[695] ;
  reg \A[696] ;
  reg \A[697] ;
  reg \A[698] ;
  reg \A[699] ;
  reg \A[7] ;
  reg \A[70] ;
  reg \A[700] ;
  reg \A[701] ;
  reg \A[702] ;
  reg \A[703] ;
  reg \A[704] ;
  reg \A[705] ;
  reg \A[706] ;
  reg \A[707] ;
  reg \A[708] ;
  reg \A[709] ;
  reg \A[71] ;
  reg \A[710] ;
  reg \A[711] ;
  reg \A[712] ;
  reg \A[713] ;
  reg \A[714] ;
  reg \A[715] ;
  reg \A[716] ;
  reg \A[717] ;
  reg \A[718] ;
  reg \A[719] ;
  reg \A[72] ;
  reg \A[720] ;
  reg \A[721] ;
  reg \A[722] ;
  reg \A[723] ;
  reg \A[724] ;
  reg \A[725] ;
  reg \A[726] ;
  reg \A[727] ;
  reg \A[728] ;
  reg \A[729] ;
  reg \A[73] ;
  reg \A[730] ;
  reg \A[731] ;
  reg \A[732] ;
  reg \A[733] ;
  reg \A[734] ;
  reg \A[735] ;
  reg \A[736] ;
  reg \A[737] ;
  reg \A[738] ;
  reg \A[739] ;
  reg \A[74] ;
  reg \A[740] ;
  reg \A[741] ;
  reg \A[742] ;
  reg \A[743] ;
  reg \A[744] ;
  reg \A[745] ;
  reg \A[746] ;
  reg \A[747] ;
  reg \A[748] ;
  reg \A[749] ;
  reg \A[75] ;
  reg \A[750] ;
  reg \A[751] ;
  reg \A[752] ;
  reg \A[753] ;
  reg \A[754] ;
  reg \A[755] ;
  reg \A[756] ;
  reg \A[757] ;
  reg \A[758] ;
  reg \A[759] ;
  reg \A[76] ;
  reg \A[760] ;
  reg \A[761] ;
  reg \A[762] ;
  reg \A[763] ;
  reg \A[764] ;
  reg \A[765] ;
  reg \A[766] ;
  reg \A[767] ;
  reg \A[768] ;
  reg \A[769] ;
  reg \A[77] ;
  reg \A[770] ;
  reg \A[771] ;
  reg \A[772] ;
  reg \A[773] ;
  reg \A[774] ;
  reg \A[775] ;
  reg \A[776] ;
  reg \A[777] ;
  reg \A[778] ;
  reg \A[779] ;
  reg \A[78] ;
  reg \A[780] ;
  reg \A[781] ;
  reg \A[782] ;
  reg \A[783] ;
  reg \A[784] ;
  reg \A[785] ;
  reg \A[786] ;
  reg \A[787] ;
  reg \A[788] ;
  reg \A[789] ;
  reg \A[79] ;
  reg \A[790] ;
  reg \A[791] ;
  reg \A[792] ;
  reg \A[793] ;
  reg \A[794] ;
  reg \A[795] ;
  reg \A[796] ;
  reg \A[797] ;
  reg \A[798] ;
  reg \A[799] ;
  reg \A[8] ;
  reg \A[80] ;
  reg \A[800] ;
  reg \A[801] ;
  reg \A[802] ;
  reg \A[803] ;
  reg \A[804] ;
  reg \A[805] ;
  reg \A[806] ;
  reg \A[807] ;
  reg \A[808] ;
  reg \A[809] ;
  reg \A[81] ;
  reg \A[810] ;
  reg \A[811] ;
  reg \A[812] ;
  reg \A[813] ;
  reg \A[814] ;
  reg \A[815] ;
  reg \A[816] ;
  reg \A[817] ;
  reg \A[818] ;
  reg \A[819] ;
  reg \A[82] ;
  reg \A[820] ;
  reg \A[821] ;
  reg \A[822] ;
  reg \A[823] ;
  reg \A[824] ;
  reg \A[825] ;
  reg \A[826] ;
  reg \A[827] ;
  reg \A[828] ;
  reg \A[829] ;
  reg \A[83] ;
  reg \A[830] ;
  reg \A[831] ;
  reg \A[832] ;
  reg \A[833] ;
  reg \A[834] ;
  reg \A[835] ;
  reg \A[836] ;
  reg \A[837] ;
  reg \A[838] ;
  reg \A[839] ;
  reg \A[84] ;
  reg \A[840] ;
  reg \A[841] ;
  reg \A[842] ;
  reg \A[843] ;
  reg \A[844] ;
  reg \A[845] ;
  reg \A[846] ;
  reg \A[847] ;
  reg \A[848] ;
  reg \A[849] ;
  reg \A[85] ;
  reg \A[850] ;
  reg \A[851] ;
  reg \A[852] ;
  reg \A[853] ;
  reg \A[854] ;
  reg \A[855] ;
  reg \A[856] ;
  reg \A[857] ;
  reg \A[858] ;
  reg \A[859] ;
  reg \A[86] ;
  reg \A[860] ;
  reg \A[861] ;
  reg \A[862] ;
  reg \A[863] ;
  reg \A[864] ;
  reg \A[865] ;
  reg \A[866] ;
  reg \A[867] ;
  reg \A[868] ;
  reg \A[869] ;
  reg \A[87] ;
  reg \A[870] ;
  reg \A[871] ;
  reg \A[872] ;
  reg \A[873] ;
  reg \A[874] ;
  reg \A[875] ;
  reg \A[876] ;
  reg \A[877] ;
  reg \A[878] ;
  reg \A[879] ;
  reg \A[88] ;
  reg \A[880] ;
  reg \A[881] ;
  reg \A[882] ;
  reg \A[883] ;
  reg \A[884] ;
  reg \A[885] ;
  reg \A[886] ;
  reg \A[887] ;
  reg \A[888] ;
  reg \A[889] ;
  reg \A[89] ;
  reg \A[890] ;
  reg \A[891] ;
  reg \A[892] ;
  reg \A[893] ;
  reg \A[894] ;
  reg \A[895] ;
  reg \A[896] ;
  reg \A[897] ;
  reg \A[898] ;
  reg \A[899] ;
  reg \A[9] ;
  reg \A[90] ;
  reg \A[900] ;
  reg \A[901] ;
  reg \A[902] ;
  reg \A[903] ;
  reg \A[904] ;
  reg \A[905] ;
  reg \A[906] ;
  reg \A[907] ;
  reg \A[908] ;
  reg \A[909] ;
  reg \A[91] ;
  reg \A[910] ;
  reg \A[911] ;
  reg \A[912] ;
  reg \A[913] ;
  reg \A[914] ;
  reg \A[915] ;
  reg \A[916] ;
  reg \A[917] ;
  reg \A[918] ;
  reg \A[919] ;
  reg \A[92] ;
  reg \A[920] ;
  reg \A[921] ;
  reg \A[922] ;
  reg \A[923] ;
  reg \A[924] ;
  reg \A[925] ;
  reg \A[926] ;
  reg \A[927] ;
  reg \A[928] ;
  reg \A[929] ;
  reg \A[93] ;
  reg \A[930] ;
  reg \A[931] ;
  reg \A[932] ;
  reg \A[933] ;
  reg \A[934] ;
  reg \A[935] ;
  reg \A[936] ;
  reg \A[937] ;
  reg \A[938] ;
  reg \A[939] ;
  reg \A[94] ;
  reg \A[940] ;
  reg \A[941] ;
  reg \A[942] ;
  reg \A[943] ;
  reg \A[944] ;
  reg \A[945] ;
  reg \A[946] ;
  reg \A[947] ;
  reg \A[948] ;
  reg \A[949] ;
  reg \A[95] ;
  reg \A[950] ;
  reg \A[951] ;
  reg \A[952] ;
  reg \A[953] ;
  reg \A[954] ;
  reg \A[955] ;
  reg \A[956] ;
  reg \A[957] ;
  reg \A[958] ;
  reg \A[959] ;
  reg \A[96] ;
  reg \A[960] ;
  reg \A[961] ;
  reg \A[962] ;
  reg \A[963] ;
  reg \A[964] ;
  reg \A[965] ;
  reg \A[966] ;
  reg \A[967] ;
  reg \A[968] ;
  reg \A[969] ;
  reg \A[97] ;
  reg \A[970] ;
  reg \A[971] ;
  reg \A[972] ;
  reg \A[973] ;
  reg \A[974] ;
  reg \A[975] ;
  reg \A[976] ;
  reg \A[977] ;
  reg \A[978] ;
  reg \A[979] ;
  reg \A[98] ;
  reg \A[980] ;
  reg \A[981] ;
  reg \A[982] ;
  reg \A[983] ;
  reg \A[984] ;
  reg \A[985] ;
  reg \A[986] ;
  reg \A[987] ;
  reg \A[988] ;
  reg \A[989] ;
  reg \A[99] ;
  reg \A[990] ;
  reg \A[991] ;
  reg \A[992] ;
  reg \A[993] ;
  reg \A[994] ;
  reg \A[995] ;
  reg \A[996] ;
  reg \A[997] ;
  reg \A[998] ;
  reg \A[999] ;
  wire maj;

  top uut (
    .\A[0] (\A[0] ),
    .\A[1] (\A[1] ),
    .\A[10] (\A[10] ),
    .\A[100] (\A[100] ),
    .\A[1000] (\A[1000] ),
    .\A[101] (\A[101] ),
    .\A[102] (\A[102] ),
    .\A[103] (\A[103] ),
    .\A[104] (\A[104] ),
    .\A[105] (\A[105] ),
    .\A[106] (\A[106] ),
    .\A[107] (\A[107] ),
    .\A[108] (\A[108] ),
    .\A[109] (\A[109] ),
    .\A[11] (\A[11] ),
    .\A[110] (\A[110] ),
    .\A[111] (\A[111] ),
    .\A[112] (\A[112] ),
    .\A[113] (\A[113] ),
    .\A[114] (\A[114] ),
    .\A[115] (\A[115] ),
    .\A[116] (\A[116] ),
    .\A[117] (\A[117] ),
    .\A[118] (\A[118] ),
    .\A[119] (\A[119] ),
    .\A[12] (\A[12] ),
    .\A[120] (\A[120] ),
    .\A[121] (\A[121] ),
    .\A[122] (\A[122] ),
    .\A[123] (\A[123] ),
    .\A[124] (\A[124] ),
    .\A[125] (\A[125] ),
    .\A[126] (\A[126] ),
    .\A[127] (\A[127] ),
    .\A[128] (\A[128] ),
    .\A[129] (\A[129] ),
    .\A[13] (\A[13] ),
    .\A[130] (\A[130] ),
    .\A[131] (\A[131] ),
    .\A[132] (\A[132] ),
    .\A[133] (\A[133] ),
    .\A[134] (\A[134] ),
    .\A[135] (\A[135] ),
    .\A[136] (\A[136] ),
    .\A[137] (\A[137] ),
    .\A[138] (\A[138] ),
    .\A[139] (\A[139] ),
    .\A[14] (\A[14] ),
    .\A[140] (\A[140] ),
    .\A[141] (\A[141] ),
    .\A[142] (\A[142] ),
    .\A[143] (\A[143] ),
    .\A[144] (\A[144] ),
    .\A[145] (\A[145] ),
    .\A[146] (\A[146] ),
    .\A[147] (\A[147] ),
    .\A[148] (\A[148] ),
    .\A[149] (\A[149] ),
    .\A[15] (\A[15] ),
    .\A[150] (\A[150] ),
    .\A[151] (\A[151] ),
    .\A[152] (\A[152] ),
    .\A[153] (\A[153] ),
    .\A[154] (\A[154] ),
    .\A[155] (\A[155] ),
    .\A[156] (\A[156] ),
    .\A[157] (\A[157] ),
    .\A[158] (\A[158] ),
    .\A[159] (\A[159] ),
    .\A[16] (\A[16] ),
    .\A[160] (\A[160] ),
    .\A[161] (\A[161] ),
    .\A[162] (\A[162] ),
    .\A[163] (\A[163] ),
    .\A[164] (\A[164] ),
    .\A[165] (\A[165] ),
    .\A[166] (\A[166] ),
    .\A[167] (\A[167] ),
    .\A[168] (\A[168] ),
    .\A[169] (\A[169] ),
    .\A[17] (\A[17] ),
    .\A[170] (\A[170] ),
    .\A[171] (\A[171] ),
    .\A[172] (\A[172] ),
    .\A[173] (\A[173] ),
    .\A[174] (\A[174] ),
    .\A[175] (\A[175] ),
    .\A[176] (\A[176] ),
    .\A[177] (\A[177] ),
    .\A[178] (\A[178] ),
    .\A[179] (\A[179] ),
    .\A[18] (\A[18] ),
    .\A[180] (\A[180] ),
    .\A[181] (\A[181] ),
    .\A[182] (\A[182] ),
    .\A[183] (\A[183] ),
    .\A[184] (\A[184] ),
    .\A[185] (\A[185] ),
    .\A[186] (\A[186] ),
    .\A[187] (\A[187] ),
    .\A[188] (\A[188] ),
    .\A[189] (\A[189] ),
    .\A[19] (\A[19] ),
    .\A[190] (\A[190] ),
    .\A[191] (\A[191] ),
    .\A[192] (\A[192] ),
    .\A[193] (\A[193] ),
    .\A[194] (\A[194] ),
    .\A[195] (\A[195] ),
    .\A[196] (\A[196] ),
    .\A[197] (\A[197] ),
    .\A[198] (\A[198] ),
    .\A[199] (\A[199] ),
    .\A[2] (\A[2] ),
    .\A[20] (\A[20] ),
    .\A[200] (\A[200] ),
    .\A[201] (\A[201] ),
    .\A[202] (\A[202] ),
    .\A[203] (\A[203] ),
    .\A[204] (\A[204] ),
    .\A[205] (\A[205] ),
    .\A[206] (\A[206] ),
    .\A[207] (\A[207] ),
    .\A[208] (\A[208] ),
    .\A[209] (\A[209] ),
    .\A[21] (\A[21] ),
    .\A[210] (\A[210] ),
    .\A[211] (\A[211] ),
    .\A[212] (\A[212] ),
    .\A[213] (\A[213] ),
    .\A[214] (\A[214] ),
    .\A[215] (\A[215] ),
    .\A[216] (\A[216] ),
    .\A[217] (\A[217] ),
    .\A[218] (\A[218] ),
    .\A[219] (\A[219] ),
    .\A[22] (\A[22] ),
    .\A[220] (\A[220] ),
    .\A[221] (\A[221] ),
    .\A[222] (\A[222] ),
    .\A[223] (\A[223] ),
    .\A[224] (\A[224] ),
    .\A[225] (\A[225] ),
    .\A[226] (\A[226] ),
    .\A[227] (\A[227] ),
    .\A[228] (\A[228] ),
    .\A[229] (\A[229] ),
    .\A[23] (\A[23] ),
    .\A[230] (\A[230] ),
    .\A[231] (\A[231] ),
    .\A[232] (\A[232] ),
    .\A[233] (\A[233] ),
    .\A[234] (\A[234] ),
    .\A[235] (\A[235] ),
    .\A[236] (\A[236] ),
    .\A[237] (\A[237] ),
    .\A[238] (\A[238] ),
    .\A[239] (\A[239] ),
    .\A[24] (\A[24] ),
    .\A[240] (\A[240] ),
    .\A[241] (\A[241] ),
    .\A[242] (\A[242] ),
    .\A[243] (\A[243] ),
    .\A[244] (\A[244] ),
    .\A[245] (\A[245] ),
    .\A[246] (\A[246] ),
    .\A[247] (\A[247] ),
    .\A[248] (\A[248] ),
    .\A[249] (\A[249] ),
    .\A[25] (\A[25] ),
    .\A[250] (\A[250] ),
    .\A[251] (\A[251] ),
    .\A[252] (\A[252] ),
    .\A[253] (\A[253] ),
    .\A[254] (\A[254] ),
    .\A[255] (\A[255] ),
    .\A[256] (\A[256] ),
    .\A[257] (\A[257] ),
    .\A[258] (\A[258] ),
    .\A[259] (\A[259] ),
    .\A[26] (\A[26] ),
    .\A[260] (\A[260] ),
    .\A[261] (\A[261] ),
    .\A[262] (\A[262] ),
    .\A[263] (\A[263] ),
    .\A[264] (\A[264] ),
    .\A[265] (\A[265] ),
    .\A[266] (\A[266] ),
    .\A[267] (\A[267] ),
    .\A[268] (\A[268] ),
    .\A[269] (\A[269] ),
    .\A[27] (\A[27] ),
    .\A[270] (\A[270] ),
    .\A[271] (\A[271] ),
    .\A[272] (\A[272] ),
    .\A[273] (\A[273] ),
    .\A[274] (\A[274] ),
    .\A[275] (\A[275] ),
    .\A[276] (\A[276] ),
    .\A[277] (\A[277] ),
    .\A[278] (\A[278] ),
    .\A[279] (\A[279] ),
    .\A[28] (\A[28] ),
    .\A[280] (\A[280] ),
    .\A[281] (\A[281] ),
    .\A[282] (\A[282] ),
    .\A[283] (\A[283] ),
    .\A[284] (\A[284] ),
    .\A[285] (\A[285] ),
    .\A[286] (\A[286] ),
    .\A[287] (\A[287] ),
    .\A[288] (\A[288] ),
    .\A[289] (\A[289] ),
    .\A[29] (\A[29] ),
    .\A[290] (\A[290] ),
    .\A[291] (\A[291] ),
    .\A[292] (\A[292] ),
    .\A[293] (\A[293] ),
    .\A[294] (\A[294] ),
    .\A[295] (\A[295] ),
    .\A[296] (\A[296] ),
    .\A[297] (\A[297] ),
    .\A[298] (\A[298] ),
    .\A[299] (\A[299] ),
    .\A[3] (\A[3] ),
    .\A[30] (\A[30] ),
    .\A[300] (\A[300] ),
    .\A[301] (\A[301] ),
    .\A[302] (\A[302] ),
    .\A[303] (\A[303] ),
    .\A[304] (\A[304] ),
    .\A[305] (\A[305] ),
    .\A[306] (\A[306] ),
    .\A[307] (\A[307] ),
    .\A[308] (\A[308] ),
    .\A[309] (\A[309] ),
    .\A[31] (\A[31] ),
    .\A[310] (\A[310] ),
    .\A[311] (\A[311] ),
    .\A[312] (\A[312] ),
    .\A[313] (\A[313] ),
    .\A[314] (\A[314] ),
    .\A[315] (\A[315] ),
    .\A[316] (\A[316] ),
    .\A[317] (\A[317] ),
    .\A[318] (\A[318] ),
    .\A[319] (\A[319] ),
    .\A[32] (\A[32] ),
    .\A[320] (\A[320] ),
    .\A[321] (\A[321] ),
    .\A[322] (\A[322] ),
    .\A[323] (\A[323] ),
    .\A[324] (\A[324] ),
    .\A[325] (\A[325] ),
    .\A[326] (\A[326] ),
    .\A[327] (\A[327] ),
    .\A[328] (\A[328] ),
    .\A[329] (\A[329] ),
    .\A[33] (\A[33] ),
    .\A[330] (\A[330] ),
    .\A[331] (\A[331] ),
    .\A[332] (\A[332] ),
    .\A[333] (\A[333] ),
    .\A[334] (\A[334] ),
    .\A[335] (\A[335] ),
    .\A[336] (\A[336] ),
    .\A[337] (\A[337] ),
    .\A[338] (\A[338] ),
    .\A[339] (\A[339] ),
    .\A[34] (\A[34] ),
    .\A[340] (\A[340] ),
    .\A[341] (\A[341] ),
    .\A[342] (\A[342] ),
    .\A[343] (\A[343] ),
    .\A[344] (\A[344] ),
    .\A[345] (\A[345] ),
    .\A[346] (\A[346] ),
    .\A[347] (\A[347] ),
    .\A[348] (\A[348] ),
    .\A[349] (\A[349] ),
    .\A[35] (\A[35] ),
    .\A[350] (\A[350] ),
    .\A[351] (\A[351] ),
    .\A[352] (\A[352] ),
    .\A[353] (\A[353] ),
    .\A[354] (\A[354] ),
    .\A[355] (\A[355] ),
    .\A[356] (\A[356] ),
    .\A[357] (\A[357] ),
    .\A[358] (\A[358] ),
    .\A[359] (\A[359] ),
    .\A[36] (\A[36] ),
    .\A[360] (\A[360] ),
    .\A[361] (\A[361] ),
    .\A[362] (\A[362] ),
    .\A[363] (\A[363] ),
    .\A[364] (\A[364] ),
    .\A[365] (\A[365] ),
    .\A[366] (\A[366] ),
    .\A[367] (\A[367] ),
    .\A[368] (\A[368] ),
    .\A[369] (\A[369] ),
    .\A[37] (\A[37] ),
    .\A[370] (\A[370] ),
    .\A[371] (\A[371] ),
    .\A[372] (\A[372] ),
    .\A[373] (\A[373] ),
    .\A[374] (\A[374] ),
    .\A[375] (\A[375] ),
    .\A[376] (\A[376] ),
    .\A[377] (\A[377] ),
    .\A[378] (\A[378] ),
    .\A[379] (\A[379] ),
    .\A[38] (\A[38] ),
    .\A[380] (\A[380] ),
    .\A[381] (\A[381] ),
    .\A[382] (\A[382] ),
    .\A[383] (\A[383] ),
    .\A[384] (\A[384] ),
    .\A[385] (\A[385] ),
    .\A[386] (\A[386] ),
    .\A[387] (\A[387] ),
    .\A[388] (\A[388] ),
    .\A[389] (\A[389] ),
    .\A[39] (\A[39] ),
    .\A[390] (\A[390] ),
    .\A[391] (\A[391] ),
    .\A[392] (\A[392] ),
    .\A[393] (\A[393] ),
    .\A[394] (\A[394] ),
    .\A[395] (\A[395] ),
    .\A[396] (\A[396] ),
    .\A[397] (\A[397] ),
    .\A[398] (\A[398] ),
    .\A[399] (\A[399] ),
    .\A[4] (\A[4] ),
    .\A[40] (\A[40] ),
    .\A[400] (\A[400] ),
    .\A[401] (\A[401] ),
    .\A[402] (\A[402] ),
    .\A[403] (\A[403] ),
    .\A[404] (\A[404] ),
    .\A[405] (\A[405] ),
    .\A[406] (\A[406] ),
    .\A[407] (\A[407] ),
    .\A[408] (\A[408] ),
    .\A[409] (\A[409] ),
    .\A[41] (\A[41] ),
    .\A[410] (\A[410] ),
    .\A[411] (\A[411] ),
    .\A[412] (\A[412] ),
    .\A[413] (\A[413] ),
    .\A[414] (\A[414] ),
    .\A[415] (\A[415] ),
    .\A[416] (\A[416] ),
    .\A[417] (\A[417] ),
    .\A[418] (\A[418] ),
    .\A[419] (\A[419] ),
    .\A[42] (\A[42] ),
    .\A[420] (\A[420] ),
    .\A[421] (\A[421] ),
    .\A[422] (\A[422] ),
    .\A[423] (\A[423] ),
    .\A[424] (\A[424] ),
    .\A[425] (\A[425] ),
    .\A[426] (\A[426] ),
    .\A[427] (\A[427] ),
    .\A[428] (\A[428] ),
    .\A[429] (\A[429] ),
    .\A[43] (\A[43] ),
    .\A[430] (\A[430] ),
    .\A[431] (\A[431] ),
    .\A[432] (\A[432] ),
    .\A[433] (\A[433] ),
    .\A[434] (\A[434] ),
    .\A[435] (\A[435] ),
    .\A[436] (\A[436] ),
    .\A[437] (\A[437] ),
    .\A[438] (\A[438] ),
    .\A[439] (\A[439] ),
    .\A[44] (\A[44] ),
    .\A[440] (\A[440] ),
    .\A[441] (\A[441] ),
    .\A[442] (\A[442] ),
    .\A[443] (\A[443] ),
    .\A[444] (\A[444] ),
    .\A[445] (\A[445] ),
    .\A[446] (\A[446] ),
    .\A[447] (\A[447] ),
    .\A[448] (\A[448] ),
    .\A[449] (\A[449] ),
    .\A[45] (\A[45] ),
    .\A[450] (\A[450] ),
    .\A[451] (\A[451] ),
    .\A[452] (\A[452] ),
    .\A[453] (\A[453] ),
    .\A[454] (\A[454] ),
    .\A[455] (\A[455] ),
    .\A[456] (\A[456] ),
    .\A[457] (\A[457] ),
    .\A[458] (\A[458] ),
    .\A[459] (\A[459] ),
    .\A[46] (\A[46] ),
    .\A[460] (\A[460] ),
    .\A[461] (\A[461] ),
    .\A[462] (\A[462] ),
    .\A[463] (\A[463] ),
    .\A[464] (\A[464] ),
    .\A[465] (\A[465] ),
    .\A[466] (\A[466] ),
    .\A[467] (\A[467] ),
    .\A[468] (\A[468] ),
    .\A[469] (\A[469] ),
    .\A[47] (\A[47] ),
    .\A[470] (\A[470] ),
    .\A[471] (\A[471] ),
    .\A[472] (\A[472] ),
    .\A[473] (\A[473] ),
    .\A[474] (\A[474] ),
    .\A[475] (\A[475] ),
    .\A[476] (\A[476] ),
    .\A[477] (\A[477] ),
    .\A[478] (\A[478] ),
    .\A[479] (\A[479] ),
    .\A[48] (\A[48] ),
    .\A[480] (\A[480] ),
    .\A[481] (\A[481] ),
    .\A[482] (\A[482] ),
    .\A[483] (\A[483] ),
    .\A[484] (\A[484] ),
    .\A[485] (\A[485] ),
    .\A[486] (\A[486] ),
    .\A[487] (\A[487] ),
    .\A[488] (\A[488] ),
    .\A[489] (\A[489] ),
    .\A[49] (\A[49] ),
    .\A[490] (\A[490] ),
    .\A[491] (\A[491] ),
    .\A[492] (\A[492] ),
    .\A[493] (\A[493] ),
    .\A[494] (\A[494] ),
    .\A[495] (\A[495] ),
    .\A[496] (\A[496] ),
    .\A[497] (\A[497] ),
    .\A[498] (\A[498] ),
    .\A[499] (\A[499] ),
    .\A[5] (\A[5] ),
    .\A[50] (\A[50] ),
    .\A[500] (\A[500] ),
    .\A[501] (\A[501] ),
    .\A[502] (\A[502] ),
    .\A[503] (\A[503] ),
    .\A[504] (\A[504] ),
    .\A[505] (\A[505] ),
    .\A[506] (\A[506] ),
    .\A[507] (\A[507] ),
    .\A[508] (\A[508] ),
    .\A[509] (\A[509] ),
    .\A[51] (\A[51] ),
    .\A[510] (\A[510] ),
    .\A[511] (\A[511] ),
    .\A[512] (\A[512] ),
    .\A[513] (\A[513] ),
    .\A[514] (\A[514] ),
    .\A[515] (\A[515] ),
    .\A[516] (\A[516] ),
    .\A[517] (\A[517] ),
    .\A[518] (\A[518] ),
    .\A[519] (\A[519] ),
    .\A[52] (\A[52] ),
    .\A[520] (\A[520] ),
    .\A[521] (\A[521] ),
    .\A[522] (\A[522] ),
    .\A[523] (\A[523] ),
    .\A[524] (\A[524] ),
    .\A[525] (\A[525] ),
    .\A[526] (\A[526] ),
    .\A[527] (\A[527] ),
    .\A[528] (\A[528] ),
    .\A[529] (\A[529] ),
    .\A[53] (\A[53] ),
    .\A[530] (\A[530] ),
    .\A[531] (\A[531] ),
    .\A[532] (\A[532] ),
    .\A[533] (\A[533] ),
    .\A[534] (\A[534] ),
    .\A[535] (\A[535] ),
    .\A[536] (\A[536] ),
    .\A[537] (\A[537] ),
    .\A[538] (\A[538] ),
    .\A[539] (\A[539] ),
    .\A[54] (\A[54] ),
    .\A[540] (\A[540] ),
    .\A[541] (\A[541] ),
    .\A[542] (\A[542] ),
    .\A[543] (\A[543] ),
    .\A[544] (\A[544] ),
    .\A[545] (\A[545] ),
    .\A[546] (\A[546] ),
    .\A[547] (\A[547] ),
    .\A[548] (\A[548] ),
    .\A[549] (\A[549] ),
    .\A[55] (\A[55] ),
    .\A[550] (\A[550] ),
    .\A[551] (\A[551] ),
    .\A[552] (\A[552] ),
    .\A[553] (\A[553] ),
    .\A[554] (\A[554] ),
    .\A[555] (\A[555] ),
    .\A[556] (\A[556] ),
    .\A[557] (\A[557] ),
    .\A[558] (\A[558] ),
    .\A[559] (\A[559] ),
    .\A[56] (\A[56] ),
    .\A[560] (\A[560] ),
    .\A[561] (\A[561] ),
    .\A[562] (\A[562] ),
    .\A[563] (\A[563] ),
    .\A[564] (\A[564] ),
    .\A[565] (\A[565] ),
    .\A[566] (\A[566] ),
    .\A[567] (\A[567] ),
    .\A[568] (\A[568] ),
    .\A[569] (\A[569] ),
    .\A[57] (\A[57] ),
    .\A[570] (\A[570] ),
    .\A[571] (\A[571] ),
    .\A[572] (\A[572] ),
    .\A[573] (\A[573] ),
    .\A[574] (\A[574] ),
    .\A[575] (\A[575] ),
    .\A[576] (\A[576] ),
    .\A[577] (\A[577] ),
    .\A[578] (\A[578] ),
    .\A[579] (\A[579] ),
    .\A[58] (\A[58] ),
    .\A[580] (\A[580] ),
    .\A[581] (\A[581] ),
    .\A[582] (\A[582] ),
    .\A[583] (\A[583] ),
    .\A[584] (\A[584] ),
    .\A[585] (\A[585] ),
    .\A[586] (\A[586] ),
    .\A[587] (\A[587] ),
    .\A[588] (\A[588] ),
    .\A[589] (\A[589] ),
    .\A[59] (\A[59] ),
    .\A[590] (\A[590] ),
    .\A[591] (\A[591] ),
    .\A[592] (\A[592] ),
    .\A[593] (\A[593] ),
    .\A[594] (\A[594] ),
    .\A[595] (\A[595] ),
    .\A[596] (\A[596] ),
    .\A[597] (\A[597] ),
    .\A[598] (\A[598] ),
    .\A[599] (\A[599] ),
    .\A[6] (\A[6] ),
    .\A[60] (\A[60] ),
    .\A[600] (\A[600] ),
    .\A[601] (\A[601] ),
    .\A[602] (\A[602] ),
    .\A[603] (\A[603] ),
    .\A[604] (\A[604] ),
    .\A[605] (\A[605] ),
    .\A[606] (\A[606] ),
    .\A[607] (\A[607] ),
    .\A[608] (\A[608] ),
    .\A[609] (\A[609] ),
    .\A[61] (\A[61] ),
    .\A[610] (\A[610] ),
    .\A[611] (\A[611] ),
    .\A[612] (\A[612] ),
    .\A[613] (\A[613] ),
    .\A[614] (\A[614] ),
    .\A[615] (\A[615] ),
    .\A[616] (\A[616] ),
    .\A[617] (\A[617] ),
    .\A[618] (\A[618] ),
    .\A[619] (\A[619] ),
    .\A[62] (\A[62] ),
    .\A[620] (\A[620] ),
    .\A[621] (\A[621] ),
    .\A[622] (\A[622] ),
    .\A[623] (\A[623] ),
    .\A[624] (\A[624] ),
    .\A[625] (\A[625] ),
    .\A[626] (\A[626] ),
    .\A[627] (\A[627] ),
    .\A[628] (\A[628] ),
    .\A[629] (\A[629] ),
    .\A[63] (\A[63] ),
    .\A[630] (\A[630] ),
    .\A[631] (\A[631] ),
    .\A[632] (\A[632] ),
    .\A[633] (\A[633] ),
    .\A[634] (\A[634] ),
    .\A[635] (\A[635] ),
    .\A[636] (\A[636] ),
    .\A[637] (\A[637] ),
    .\A[638] (\A[638] ),
    .\A[639] (\A[639] ),
    .\A[64] (\A[64] ),
    .\A[640] (\A[640] ),
    .\A[641] (\A[641] ),
    .\A[642] (\A[642] ),
    .\A[643] (\A[643] ),
    .\A[644] (\A[644] ),
    .\A[645] (\A[645] ),
    .\A[646] (\A[646] ),
    .\A[647] (\A[647] ),
    .\A[648] (\A[648] ),
    .\A[649] (\A[649] ),
    .\A[65] (\A[65] ),
    .\A[650] (\A[650] ),
    .\A[651] (\A[651] ),
    .\A[652] (\A[652] ),
    .\A[653] (\A[653] ),
    .\A[654] (\A[654] ),
    .\A[655] (\A[655] ),
    .\A[656] (\A[656] ),
    .\A[657] (\A[657] ),
    .\A[658] (\A[658] ),
    .\A[659] (\A[659] ),
    .\A[66] (\A[66] ),
    .\A[660] (\A[660] ),
    .\A[661] (\A[661] ),
    .\A[662] (\A[662] ),
    .\A[663] (\A[663] ),
    .\A[664] (\A[664] ),
    .\A[665] (\A[665] ),
    .\A[666] (\A[666] ),
    .\A[667] (\A[667] ),
    .\A[668] (\A[668] ),
    .\A[669] (\A[669] ),
    .\A[67] (\A[67] ),
    .\A[670] (\A[670] ),
    .\A[671] (\A[671] ),
    .\A[672] (\A[672] ),
    .\A[673] (\A[673] ),
    .\A[674] (\A[674] ),
    .\A[675] (\A[675] ),
    .\A[676] (\A[676] ),
    .\A[677] (\A[677] ),
    .\A[678] (\A[678] ),
    .\A[679] (\A[679] ),
    .\A[68] (\A[68] ),
    .\A[680] (\A[680] ),
    .\A[681] (\A[681] ),
    .\A[682] (\A[682] ),
    .\A[683] (\A[683] ),
    .\A[684] (\A[684] ),
    .\A[685] (\A[685] ),
    .\A[686] (\A[686] ),
    .\A[687] (\A[687] ),
    .\A[688] (\A[688] ),
    .\A[689] (\A[689] ),
    .\A[69] (\A[69] ),
    .\A[690] (\A[690] ),
    .\A[691] (\A[691] ),
    .\A[692] (\A[692] ),
    .\A[693] (\A[693] ),
    .\A[694] (\A[694] ),
    .\A[695] (\A[695] ),
    .\A[696] (\A[696] ),
    .\A[697] (\A[697] ),
    .\A[698] (\A[698] ),
    .\A[699] (\A[699] ),
    .\A[7] (\A[7] ),
    .\A[70] (\A[70] ),
    .\A[700] (\A[700] ),
    .\A[701] (\A[701] ),
    .\A[702] (\A[702] ),
    .\A[703] (\A[703] ),
    .\A[704] (\A[704] ),
    .\A[705] (\A[705] ),
    .\A[706] (\A[706] ),
    .\A[707] (\A[707] ),
    .\A[708] (\A[708] ),
    .\A[709] (\A[709] ),
    .\A[71] (\A[71] ),
    .\A[710] (\A[710] ),
    .\A[711] (\A[711] ),
    .\A[712] (\A[712] ),
    .\A[713] (\A[713] ),
    .\A[714] (\A[714] ),
    .\A[715] (\A[715] ),
    .\A[716] (\A[716] ),
    .\A[717] (\A[717] ),
    .\A[718] (\A[718] ),
    .\A[719] (\A[719] ),
    .\A[72] (\A[72] ),
    .\A[720] (\A[720] ),
    .\A[721] (\A[721] ),
    .\A[722] (\A[722] ),
    .\A[723] (\A[723] ),
    .\A[724] (\A[724] ),
    .\A[725] (\A[725] ),
    .\A[726] (\A[726] ),
    .\A[727] (\A[727] ),
    .\A[728] (\A[728] ),
    .\A[729] (\A[729] ),
    .\A[73] (\A[73] ),
    .\A[730] (\A[730] ),
    .\A[731] (\A[731] ),
    .\A[732] (\A[732] ),
    .\A[733] (\A[733] ),
    .\A[734] (\A[734] ),
    .\A[735] (\A[735] ),
    .\A[736] (\A[736] ),
    .\A[737] (\A[737] ),
    .\A[738] (\A[738] ),
    .\A[739] (\A[739] ),
    .\A[74] (\A[74] ),
    .\A[740] (\A[740] ),
    .\A[741] (\A[741] ),
    .\A[742] (\A[742] ),
    .\A[743] (\A[743] ),
    .\A[744] (\A[744] ),
    .\A[745] (\A[745] ),
    .\A[746] (\A[746] ),
    .\A[747] (\A[747] ),
    .\A[748] (\A[748] ),
    .\A[749] (\A[749] ),
    .\A[75] (\A[75] ),
    .\A[750] (\A[750] ),
    .\A[751] (\A[751] ),
    .\A[752] (\A[752] ),
    .\A[753] (\A[753] ),
    .\A[754] (\A[754] ),
    .\A[755] (\A[755] ),
    .\A[756] (\A[756] ),
    .\A[757] (\A[757] ),
    .\A[758] (\A[758] ),
    .\A[759] (\A[759] ),
    .\A[76] (\A[76] ),
    .\A[760] (\A[760] ),
    .\A[761] (\A[761] ),
    .\A[762] (\A[762] ),
    .\A[763] (\A[763] ),
    .\A[764] (\A[764] ),
    .\A[765] (\A[765] ),
    .\A[766] (\A[766] ),
    .\A[767] (\A[767] ),
    .\A[768] (\A[768] ),
    .\A[769] (\A[769] ),
    .\A[77] (\A[77] ),
    .\A[770] (\A[770] ),
    .\A[771] (\A[771] ),
    .\A[772] (\A[772] ),
    .\A[773] (\A[773] ),
    .\A[774] (\A[774] ),
    .\A[775] (\A[775] ),
    .\A[776] (\A[776] ),
    .\A[777] (\A[777] ),
    .\A[778] (\A[778] ),
    .\A[779] (\A[779] ),
    .\A[78] (\A[78] ),
    .\A[780] (\A[780] ),
    .\A[781] (\A[781] ),
    .\A[782] (\A[782] ),
    .\A[783] (\A[783] ),
    .\A[784] (\A[784] ),
    .\A[785] (\A[785] ),
    .\A[786] (\A[786] ),
    .\A[787] (\A[787] ),
    .\A[788] (\A[788] ),
    .\A[789] (\A[789] ),
    .\A[79] (\A[79] ),
    .\A[790] (\A[790] ),
    .\A[791] (\A[791] ),
    .\A[792] (\A[792] ),
    .\A[793] (\A[793] ),
    .\A[794] (\A[794] ),
    .\A[795] (\A[795] ),
    .\A[796] (\A[796] ),
    .\A[797] (\A[797] ),
    .\A[798] (\A[798] ),
    .\A[799] (\A[799] ),
    .\A[8] (\A[8] ),
    .\A[80] (\A[80] ),
    .\A[800] (\A[800] ),
    .\A[801] (\A[801] ),
    .\A[802] (\A[802] ),
    .\A[803] (\A[803] ),
    .\A[804] (\A[804] ),
    .\A[805] (\A[805] ),
    .\A[806] (\A[806] ),
    .\A[807] (\A[807] ),
    .\A[808] (\A[808] ),
    .\A[809] (\A[809] ),
    .\A[81] (\A[81] ),
    .\A[810] (\A[810] ),
    .\A[811] (\A[811] ),
    .\A[812] (\A[812] ),
    .\A[813] (\A[813] ),
    .\A[814] (\A[814] ),
    .\A[815] (\A[815] ),
    .\A[816] (\A[816] ),
    .\A[817] (\A[817] ),
    .\A[818] (\A[818] ),
    .\A[819] (\A[819] ),
    .\A[82] (\A[82] ),
    .\A[820] (\A[820] ),
    .\A[821] (\A[821] ),
    .\A[822] (\A[822] ),
    .\A[823] (\A[823] ),
    .\A[824] (\A[824] ),
    .\A[825] (\A[825] ),
    .\A[826] (\A[826] ),
    .\A[827] (\A[827] ),
    .\A[828] (\A[828] ),
    .\A[829] (\A[829] ),
    .\A[83] (\A[83] ),
    .\A[830] (\A[830] ),
    .\A[831] (\A[831] ),
    .\A[832] (\A[832] ),
    .\A[833] (\A[833] ),
    .\A[834] (\A[834] ),
    .\A[835] (\A[835] ),
    .\A[836] (\A[836] ),
    .\A[837] (\A[837] ),
    .\A[838] (\A[838] ),
    .\A[839] (\A[839] ),
    .\A[84] (\A[84] ),
    .\A[840] (\A[840] ),
    .\A[841] (\A[841] ),
    .\A[842] (\A[842] ),
    .\A[843] (\A[843] ),
    .\A[844] (\A[844] ),
    .\A[845] (\A[845] ),
    .\A[846] (\A[846] ),
    .\A[847] (\A[847] ),
    .\A[848] (\A[848] ),
    .\A[849] (\A[849] ),
    .\A[85] (\A[85] ),
    .\A[850] (\A[850] ),
    .\A[851] (\A[851] ),
    .\A[852] (\A[852] ),
    .\A[853] (\A[853] ),
    .\A[854] (\A[854] ),
    .\A[855] (\A[855] ),
    .\A[856] (\A[856] ),
    .\A[857] (\A[857] ),
    .\A[858] (\A[858] ),
    .\A[859] (\A[859] ),
    .\A[86] (\A[86] ),
    .\A[860] (\A[860] ),
    .\A[861] (\A[861] ),
    .\A[862] (\A[862] ),
    .\A[863] (\A[863] ),
    .\A[864] (\A[864] ),
    .\A[865] (\A[865] ),
    .\A[866] (\A[866] ),
    .\A[867] (\A[867] ),
    .\A[868] (\A[868] ),
    .\A[869] (\A[869] ),
    .\A[87] (\A[87] ),
    .\A[870] (\A[870] ),
    .\A[871] (\A[871] ),
    .\A[872] (\A[872] ),
    .\A[873] (\A[873] ),
    .\A[874] (\A[874] ),
    .\A[875] (\A[875] ),
    .\A[876] (\A[876] ),
    .\A[877] (\A[877] ),
    .\A[878] (\A[878] ),
    .\A[879] (\A[879] ),
    .\A[88] (\A[88] ),
    .\A[880] (\A[880] ),
    .\A[881] (\A[881] ),
    .\A[882] (\A[882] ),
    .\A[883] (\A[883] ),
    .\A[884] (\A[884] ),
    .\A[885] (\A[885] ),
    .\A[886] (\A[886] ),
    .\A[887] (\A[887] ),
    .\A[888] (\A[888] ),
    .\A[889] (\A[889] ),
    .\A[89] (\A[89] ),
    .\A[890] (\A[890] ),
    .\A[891] (\A[891] ),
    .\A[892] (\A[892] ),
    .\A[893] (\A[893] ),
    .\A[894] (\A[894] ),
    .\A[895] (\A[895] ),
    .\A[896] (\A[896] ),
    .\A[897] (\A[897] ),
    .\A[898] (\A[898] ),
    .\A[899] (\A[899] ),
    .\A[9] (\A[9] ),
    .\A[90] (\A[90] ),
    .\A[900] (\A[900] ),
    .\A[901] (\A[901] ),
    .\A[902] (\A[902] ),
    .\A[903] (\A[903] ),
    .\A[904] (\A[904] ),
    .\A[905] (\A[905] ),
    .\A[906] (\A[906] ),
    .\A[907] (\A[907] ),
    .\A[908] (\A[908] ),
    .\A[909] (\A[909] ),
    .\A[91] (\A[91] ),
    .\A[910] (\A[910] ),
    .\A[911] (\A[911] ),
    .\A[912] (\A[912] ),
    .\A[913] (\A[913] ),
    .\A[914] (\A[914] ),
    .\A[915] (\A[915] ),
    .\A[916] (\A[916] ),
    .\A[917] (\A[917] ),
    .\A[918] (\A[918] ),
    .\A[919] (\A[919] ),
    .\A[92] (\A[92] ),
    .\A[920] (\A[920] ),
    .\A[921] (\A[921] ),
    .\A[922] (\A[922] ),
    .\A[923] (\A[923] ),
    .\A[924] (\A[924] ),
    .\A[925] (\A[925] ),
    .\A[926] (\A[926] ),
    .\A[927] (\A[927] ),
    .\A[928] (\A[928] ),
    .\A[929] (\A[929] ),
    .\A[93] (\A[93] ),
    .\A[930] (\A[930] ),
    .\A[931] (\A[931] ),
    .\A[932] (\A[932] ),
    .\A[933] (\A[933] ),
    .\A[934] (\A[934] ),
    .\A[935] (\A[935] ),
    .\A[936] (\A[936] ),
    .\A[937] (\A[937] ),
    .\A[938] (\A[938] ),
    .\A[939] (\A[939] ),
    .\A[94] (\A[94] ),
    .\A[940] (\A[940] ),
    .\A[941] (\A[941] ),
    .\A[942] (\A[942] ),
    .\A[943] (\A[943] ),
    .\A[944] (\A[944] ),
    .\A[945] (\A[945] ),
    .\A[946] (\A[946] ),
    .\A[947] (\A[947] ),
    .\A[948] (\A[948] ),
    .\A[949] (\A[949] ),
    .\A[95] (\A[95] ),
    .\A[950] (\A[950] ),
    .\A[951] (\A[951] ),
    .\A[952] (\A[952] ),
    .\A[953] (\A[953] ),
    .\A[954] (\A[954] ),
    .\A[955] (\A[955] ),
    .\A[956] (\A[956] ),
    .\A[957] (\A[957] ),
    .\A[958] (\A[958] ),
    .\A[959] (\A[959] ),
    .\A[96] (\A[96] ),
    .\A[960] (\A[960] ),
    .\A[961] (\A[961] ),
    .\A[962] (\A[962] ),
    .\A[963] (\A[963] ),
    .\A[964] (\A[964] ),
    .\A[965] (\A[965] ),
    .\A[966] (\A[966] ),
    .\A[967] (\A[967] ),
    .\A[968] (\A[968] ),
    .\A[969] (\A[969] ),
    .\A[97] (\A[97] ),
    .\A[970] (\A[970] ),
    .\A[971] (\A[971] ),
    .\A[972] (\A[972] ),
    .\A[973] (\A[973] ),
    .\A[974] (\A[974] ),
    .\A[975] (\A[975] ),
    .\A[976] (\A[976] ),
    .\A[977] (\A[977] ),
    .\A[978] (\A[978] ),
    .\A[979] (\A[979] ),
    .\A[98] (\A[98] ),
    .\A[980] (\A[980] ),
    .\A[981] (\A[981] ),
    .\A[982] (\A[982] ),
    .\A[983] (\A[983] ),
    .\A[984] (\A[984] ),
    .\A[985] (\A[985] ),
    .\A[986] (\A[986] ),
    .\A[987] (\A[987] ),
    .\A[988] (\A[988] ),
    .\A[989] (\A[989] ),
    .\A[99] (\A[99] ),
    .\A[990] (\A[990] ),
    .\A[991] (\A[991] ),
    .\A[992] (\A[992] ),
    .\A[993] (\A[993] ),
    .\A[994] (\A[994] ),
    .\A[995] (\A[995] ),
    .\A[996] (\A[996] ),
    .\A[997] (\A[997] ),
    .\A[998] (\A[998] ),
    .\A[999] (\A[999] ),
    .maj (maj)
  );

  integer i;
  parameter STEPS = 2048;
  parameter PRINT_EVERY = 16;

  initial begin
    // 初始化: V16策略 - 精细选择性探测
    \A[0] = 1'b0;
    \A[1] = 1'b0;
    \A[2] = 1'b0;
    \A[3] = 1'b0;
    \A[4] = 1'b0;
    \A[5] = 1'b0;
    \A[6] = 1'b0;
    \A[7] = 1'b0;
    \A[8] = 1'b0;
    \A[9] = 1'b0;
    \A[10] = 1'b0;
    \A[11] = 1'b0;
    \A[12] = 1'b0;
    \A[13] = 1'b0;
    \A[14] = 1'b0;
    \A[15] = 1'b0;
    \A[16] = 1'b0;
    \A[17] = 1'b0;
    \A[18] = 1'b0;
    \A[19] = 1'b0;
    \A[20] = 1'b0;
    \A[21] = 1'b0;
    \A[22] = 1'b0;
    \A[23] = 1'b0;
    \A[24] = 1'b0;
    \A[25] = 1'b0;
    \A[26] = 1'b0;
    \A[27] = 1'b0;
    \A[28] = 1'b0;
    \A[29] = 1'b0;
    \A[30] = 1'b0;
    \A[31] = 1'b0;
    \A[32] = 1'b0;
    \A[33] = 1'b0;
    \A[34] = 1'b0;
    \A[35] = 1'b0;
    \A[36] = 1'b0;
    \A[37] = 1'b0;
    \A[38] = 1'b0;
    \A[39] = 1'b0;
    \A[40] = 1'b0;
    \A[41] = 1'b0;
    \A[42] = 1'b0;
    \A[43] = 1'b0;
    \A[44] = 1'b0;
    \A[45] = 1'b0;
    \A[46] = 1'b0;
    \A[47] = 1'b0;
    \A[48] = 1'b0;
    \A[49] = 1'b0;
    \A[50] = 1'b0;
    \A[51] = 1'b0;
    \A[52] = 1'b0;
    \A[53] = 1'b0;
    \A[54] = 1'b0;
    \A[55] = 1'b0;
    \A[56] = 1'b0;
    \A[57] = 1'b0;
    \A[58] = 1'b0;
    \A[59] = 1'b0;
    \A[60] = 1'b0;
    \A[61] = 1'b0;
    \A[62] = 1'b0;
    \A[63] = 1'b0;
    \A[64] = 1'b1;
    \A[65] = 1'b1;
    \A[66] = 1'b1;
    \A[67] = 1'b1;
    \A[68] = 1'b1;
    \A[69] = 1'b1;
    \A[70] = 1'b1;
    \A[71] = 1'b1;
    \A[72] = 1'b1;
    \A[73] = 1'b1;
    \A[74] = 1'b1;
    \A[75] = 1'b1;
    \A[76] = 1'b1;
    \A[77] = 1'b1;
    \A[78] = 1'b1;
    \A[79] = 1'b1;
    \A[80] = 1'b1;
    \A[81] = 1'b1;
    \A[82] = 1'b1;
    \A[83] = 1'b1;
    \A[84] = 1'b1;
    \A[85] = 1'b1;
    \A[86] = 1'b1;
    \A[87] = 1'b1;
    \A[88] = 1'b1;
    \A[89] = 1'b1;
    \A[90] = 1'b1;
    \A[91] = 1'b1;
    \A[92] = 1'b1;
    \A[93] = 1'b1;
    \A[94] = 1'b1;
    \A[95] = 1'b1;
    \A[96] = 1'b1;
    \A[97] = 1'b1;
    \A[98] = 1'b1;
    \A[99] = 1'b1;
    \A[100] = 1'b1;
    \A[101] = 1'b1;
    \A[102] = 1'b1;
    \A[103] = 1'b1;
    \A[104] = 1'b1;
    \A[105] = 1'b1;
    \A[106] = 1'b1;
    \A[107] = 1'b1;
    \A[108] = 1'b1;
    \A[109] = 1'b1;
    \A[110] = 1'b1;
    \A[111] = 1'b1;
    \A[112] = 1'b1;
    \A[113] = 1'b1;
    \A[114] = 1'b1;
    \A[115] = 1'b1;
    \A[116] = 1'b1;
    \A[117] = 1'b1;
    \A[118] = 1'b1;
    \A[119] = 1'b1;
    \A[120] = 1'b1;
    \A[121] = 1'b1;
    \A[122] = 1'b1;
    \A[123] = 1'b1;
    \A[124] = 1'b1;
    \A[125] = 1'b1;
    \A[126] = 1'b1;
    \A[127] = 1'b1;
    \A[128] = 1'b1;
    \A[129] = 1'b1;
    \A[130] = 1'b1;
    \A[131] = 1'b1;
    \A[132] = 1'b1;
    \A[133] = 1'b1;
    \A[134] = 1'b1;
    \A[135] = 1'b1;
    \A[136] = 1'b1;
    \A[137] = 1'b1;
    \A[138] = 1'b1;
    \A[139] = 1'b1;
    \A[140] = 1'b1;
    \A[141] = 1'b1;
    \A[142] = 1'b1;
    \A[143] = 1'b1;
    \A[144] = 1'b1;
    \A[145] = 1'b1;
    \A[146] = 1'b1;
    \A[147] = 1'b1;
    \A[148] = 1'b1;
    \A[149] = 1'b1;
    \A[150] = 1'b1;
    \A[151] = 1'b1;
    \A[152] = 1'b1;
    \A[153] = 1'b1;
    \A[154] = 1'b1;
    \A[155] = 1'b1;
    \A[156] = 1'b1;
    \A[157] = 1'b1;
    \A[158] = 1'b1;
    \A[159] = 1'b1;
    \A[160] = 1'b1;
    \A[161] = 1'b1;
    \A[162] = 1'b1;
    \A[163] = 1'b1;
    \A[164] = 1'b1;
    \A[165] = 1'b1;
    \A[166] = 1'b1;
    \A[167] = 1'b1;
    \A[168] = 1'b1;
    \A[169] = 1'b1;
    \A[170] = 1'b1;
    \A[171] = 1'b1;
    \A[172] = 1'b1;
    \A[173] = 1'b1;
    \A[174] = 1'b1;
    \A[175] = 1'b1;
    \A[176] = 1'b1;
    \A[177] = 1'b1;
    \A[178] = 1'b1;
    \A[179] = 1'b1;
    \A[180] = 1'b1;
    \A[181] = 1'b1;
    \A[182] = 1'b1;
    \A[183] = 1'b1;
    \A[184] = 1'b1;
    \A[185] = 1'b1;
    \A[186] = 1'b1;
    \A[187] = 1'b1;
    \A[188] = 1'b1;
    \A[189] = 1'b1;
    \A[190] = 1'b1;
    \A[191] = 1'b1;
    \A[192] = 1'b1;
    \A[193] = 1'b1;
    \A[194] = 1'b1;
    \A[195] = 1'b1;
    \A[196] = 1'b1;
    \A[197] = 1'b1;
    \A[198] = 1'b1;
    \A[199] = 1'b1;
    \A[200] = 1'b1;
    \A[201] = 1'b1;
    \A[202] = 1'b1;
    \A[203] = 1'b1;
    \A[204] = 1'b1;
    \A[205] = 1'b1;
    \A[206] = 1'b1;
    \A[207] = 1'b1;
    \A[208] = 1'b1;
    \A[209] = 1'b1;
    \A[210] = 1'b1;
    \A[211] = 1'b1;
    \A[212] = 1'b1;
    \A[213] = 1'b1;
    \A[214] = 1'b1;
    \A[215] = 1'b1;
    \A[216] = 1'b1;
    \A[217] = 1'b1;
    \A[218] = 1'b1;
    \A[219] = 1'b1;
    \A[220] = 1'b1;
    \A[221] = 1'b1;
    \A[222] = 1'b1;
    \A[223] = 1'b1;
    \A[224] = 1'b1;
    \A[225] = 1'b1;
    \A[226] = 1'b1;
    \A[227] = 1'b1;
    \A[228] = 1'b1;
    \A[229] = 1'b1;
    \A[230] = 1'b1;
    \A[231] = 1'b1;
    \A[232] = 1'b1;
    \A[233] = 1'b1;
    \A[234] = 1'b1;
    \A[235] = 1'b1;
    \A[236] = 1'b1;
    \A[237] = 1'b1;
    \A[238] = 1'b1;
    \A[239] = 1'b1;
    \A[240] = 1'b1;
    \A[241] = 1'b1;
    \A[242] = 1'b1;
    \A[243] = 1'b1;
    \A[244] = 1'b1;
    \A[245] = 1'b1;
    \A[246] = 1'b1;
    \A[247] = 1'b1;
    \A[248] = 1'b1;
    \A[249] = 1'b1;
    \A[250] = 1'b1;
    \A[251] = 1'b1;
    \A[252] = 1'b1;
    \A[253] = 1'b1;
    \A[254] = 1'b1;
    \A[255] = 1'b1;
    \A[256] = 1'b1;
    \A[257] = 1'b1;
    \A[258] = 1'b1;
    \A[259] = 1'b1;
    \A[260] = 1'b1;
    \A[261] = 1'b1;
    \A[262] = 1'b1;
    \A[263] = 1'b1;
    \A[264] = 1'b1;
    \A[265] = 1'b1;
    \A[266] = 1'b1;
    \A[267] = 1'b1;
    \A[268] = 1'b1;
    \A[269] = 1'b1;
    \A[270] = 1'b1;
    \A[271] = 1'b1;
    \A[272] = 1'b1;
    \A[273] = 1'b1;
    \A[274] = 1'b1;
    \A[275] = 1'b1;
    \A[276] = 1'b1;
    \A[277] = 1'b1;
    \A[278] = 1'b1;
    \A[279] = 1'b1;
    \A[280] = 1'b1;
    \A[281] = 1'b1;
    \A[282] = 1'b1;
    \A[283] = 1'b1;
    \A[284] = 1'b1;
    \A[285] = 1'b1;
    \A[286] = 1'b1;
    \A[287] = 1'b1;
    \A[288] = 1'b1;
    \A[289] = 1'b1;
    \A[290] = 1'b1;
    \A[291] = 1'b1;
    \A[292] = 1'b1;
    \A[293] = 1'b1;
    \A[294] = 1'b1;
    \A[295] = 1'b1;
    \A[296] = 1'b1;
    \A[297] = 1'b1;
    \A[298] = 1'b1;
    \A[299] = 1'b1;
    \A[300] = 1'b1;
    \A[301] = 1'b1;
    \A[302] = 1'b1;
    \A[303] = 1'b1;
    \A[304] = 1'b1;
    \A[305] = 1'b1;
    \A[306] = 1'b1;
    \A[307] = 1'b1;
    \A[308] = 1'b1;
    \A[309] = 1'b1;
    \A[310] = 1'b1;
    \A[311] = 1'b1;
    \A[312] = 1'b1;
    \A[313] = 1'b1;
    \A[314] = 1'b1;
    \A[315] = 1'b1;
    \A[316] = 1'b1;
    \A[317] = 1'b1;
    \A[318] = 1'b1;
    \A[319] = 1'b1;
    \A[320] = 1'b1;
    \A[321] = 1'b1;
    \A[322] = 1'b1;
    \A[323] = 1'b1;
    \A[324] = 1'b1;
    \A[325] = 1'b1;
    \A[326] = 1'b1;
    \A[327] = 1'b1;
    \A[328] = 1'b1;
    \A[329] = 1'b1;
    \A[330] = 1'b1;
    \A[331] = 1'b1;
    \A[332] = 1'b1;
    \A[333] = 1'b1;
    \A[334] = 1'b1;
    \A[335] = 1'b1;
    \A[336] = 1'b1;
    \A[337] = 1'b1;
    \A[338] = 1'b1;
    \A[339] = 1'b1;
    \A[340] = 1'b1;
    \A[341] = 1'b1;
    \A[342] = 1'b1;
    \A[343] = 1'b1;
    \A[344] = 1'b1;
    \A[345] = 1'b1;
    \A[346] = 1'b1;
    \A[347] = 1'b1;
    \A[348] = 1'b1;
    \A[349] = 1'b1;
    \A[350] = 1'b1;
    \A[351] = 1'b1;
    \A[352] = 1'b1;
    \A[353] = 1'b1;
    \A[354] = 1'b1;
    \A[355] = 1'b1;
    \A[356] = 1'b1;
    \A[357] = 1'b1;
    \A[358] = 1'b1;
    \A[359] = 1'b1;
    \A[360] = 1'b1;
    \A[361] = 1'b1;
    \A[362] = 1'b1;
    \A[363] = 1'b1;
    \A[364] = 1'b1;
    \A[365] = 1'b1;
    \A[366] = 1'b1;
    \A[367] = 1'b1;
    \A[368] = 1'b1;
    \A[369] = 1'b1;
    \A[370] = 1'b1;
    \A[371] = 1'b1;
    \A[372] = 1'b1;
    \A[373] = 1'b1;
    \A[374] = 1'b1;
    \A[375] = 1'b1;
    \A[376] = 1'b1;
    \A[377] = 1'b1;
    \A[378] = 1'b1;
    \A[379] = 1'b1;
    \A[380] = 1'b1;
    \A[381] = 1'b1;
    \A[382] = 1'b1;
    \A[383] = 1'b1;
    \A[384] = 1'b1;
    \A[385] = 1'b1;
    \A[386] = 1'b1;
    \A[387] = 1'b1;
    \A[388] = 1'b1;
    \A[389] = 1'b1;
    \A[390] = 1'b1;
    \A[391] = 1'b1;
    \A[392] = 1'b1;
    \A[393] = 1'b1;
    \A[394] = 1'b1;
    \A[395] = 1'b1;
    \A[396] = 1'b1;
    \A[397] = 1'b1;
    \A[398] = 1'b1;
    \A[399] = 1'b1;
    \A[400] = 1'b1;
    \A[401] = 1'b1;
    \A[402] = 1'b1;
    \A[403] = 1'b1;
    \A[404] = 1'b1;
    \A[405] = 1'b1;
    \A[406] = 1'b1;
    \A[407] = 1'b1;
    \A[408] = 1'b1;
    \A[409] = 1'b1;
    \A[410] = 1'b1;
    \A[411] = 1'b1;
    \A[412] = 1'b1;
    \A[413] = 1'b1;
    \A[414] = 1'b1;
    \A[415] = 1'b1;
    \A[416] = 1'b1;
    \A[417] = 1'b1;
    \A[418] = 1'b1;
    \A[419] = 1'b1;
    \A[420] = 1'b1;
    \A[421] = 1'b1;
    \A[422] = 1'b1;
    \A[423] = 1'b1;
    \A[424] = 1'b1;
    \A[425] = 1'b1;
    \A[426] = 1'b1;
    \A[427] = 1'b1;
    \A[428] = 1'b1;
    \A[429] = 1'b1;
    \A[430] = 1'b1;
    \A[431] = 1'b1;
    \A[432] = 1'b1;
    \A[433] = 1'b1;
    \A[434] = 1'b1;
    \A[435] = 1'b1;
    \A[436] = 1'b1;
    \A[437] = 1'b1;
    \A[438] = 1'b1;
    \A[439] = 1'b1;
    \A[440] = 1'b1;
    \A[441] = 1'b1;
    \A[442] = 1'b1;
    \A[443] = 1'b1;
    \A[444] = 1'b1;
    \A[445] = 1'b1;
    \A[446] = 1'b1;
    \A[447] = 1'b1;
    \A[448] = 1'b1;
    \A[449] = 1'b1;
    \A[450] = 1'b1;
    \A[451] = 1'b1;
    \A[452] = 1'b1;
    \A[453] = 1'b1;
    \A[454] = 1'b1;
    \A[455] = 1'b1;
    \A[456] = 1'b1;
    \A[457] = 1'b1;
    \A[458] = 1'b1;
    \A[459] = 1'b1;
    \A[460] = 1'b1;
    \A[461] = 1'b1;
    \A[462] = 1'b1;
    \A[463] = 1'b1;
    \A[464] = 1'b1;
    \A[465] = 1'b1;
    \A[466] = 1'b1;
    \A[467] = 1'b1;
    \A[468] = 1'b1;
    \A[469] = 1'b1;
    \A[470] = 1'b1;
    \A[471] = 1'b1;
    \A[472] = 1'b1;
    \A[473] = 1'b1;
    \A[474] = 1'b1;
    \A[475] = 1'b1;
    \A[476] = 1'b1;
    \A[477] = 1'b1;
    \A[478] = 1'b1;
    \A[479] = 1'b1;
    \A[480] = 1'b1;
    \A[481] = 1'b1;
    \A[482] = 1'b1;
    \A[483] = 1'b1;
    \A[484] = 1'b1;
    \A[485] = 1'b1;
    \A[486] = 1'b1;
    \A[487] = 1'b1;
    \A[488] = 1'b1;
    \A[489] = 1'b1;
    \A[490] = 1'b1;
    \A[491] = 1'b1;
    \A[492] = 1'b1;
    \A[493] = 1'b1;
    \A[494] = 1'b1;
    \A[495] = 1'b1;
    \A[496] = 1'b1;
    \A[497] = 1'b1;
    \A[498] = 1'b1;
    \A[499] = 1'b0;
    \A[500] = 1'b0;
    \A[501] = 1'b0;
    \A[502] = 1'b0;
    \A[503] = 1'b0;
    \A[504] = 1'b0;
    \A[505] = 1'b0;
    \A[506] = 1'b0;
    \A[507] = 1'b0;
    \A[508] = 1'b0;
    \A[509] = 1'b0;
    \A[510] = 1'b0;
    \A[511] = 1'b0;
    \A[512] = 1'b0;
    \A[513] = 1'b0;
    \A[514] = 1'b0;
    \A[515] = 1'b0;
    \A[516] = 1'b0;
    \A[517] = 1'b0;
    \A[518] = 1'b0;
    \A[519] = 1'b0;
    \A[520] = 1'b0;
    \A[521] = 1'b0;
    \A[522] = 1'b0;
    \A[523] = 1'b0;
    \A[524] = 1'b0;
    \A[525] = 1'b0;
    \A[526] = 1'b0;
    \A[527] = 1'b0;
    \A[528] = 1'b0;
    \A[529] = 1'b0;
    \A[530] = 1'b0;
    \A[531] = 1'b0;
    \A[532] = 1'b0;
    \A[533] = 1'b0;
    \A[534] = 1'b0;
    \A[535] = 1'b0;
    \A[536] = 1'b0;
    \A[537] = 1'b0;
    \A[538] = 1'b0;
    \A[539] = 1'b0;
    \A[540] = 1'b0;
    \A[541] = 1'b0;
    \A[542] = 1'b0;
    \A[543] = 1'b0;
    \A[544] = 1'b0;
    \A[545] = 1'b0;
    \A[546] = 1'b0;
    \A[547] = 1'b0;
    \A[548] = 1'b0;
    \A[549] = 1'b0;
    \A[550] = 1'b0;
    \A[551] = 1'b0;
    \A[552] = 1'b0;
    \A[553] = 1'b0;
    \A[554] = 1'b0;
    \A[555] = 1'b0;
    \A[556] = 1'b0;
    \A[557] = 1'b0;
    \A[558] = 1'b0;
    \A[559] = 1'b0;
    \A[560] = 1'b0;
    \A[561] = 1'b0;
    \A[562] = 1'b0;
    \A[563] = 1'b0;
    \A[564] = 1'b0;
    \A[565] = 1'b0;
    \A[566] = 1'b0;
    \A[567] = 1'b0;
    \A[568] = 1'b0;
    \A[569] = 1'b0;
    \A[570] = 1'b0;
    \A[571] = 1'b0;
    \A[572] = 1'b0;
    \A[573] = 1'b0;
    \A[574] = 1'b0;
    \A[575] = 1'b0;
    \A[576] = 1'b0;
    \A[577] = 1'b0;
    \A[578] = 1'b0;
    \A[579] = 1'b0;
    \A[580] = 1'b0;
    \A[581] = 1'b0;
    \A[582] = 1'b0;
    \A[583] = 1'b0;
    \A[584] = 1'b0;
    \A[585] = 1'b0;
    \A[586] = 1'b0;
    \A[587] = 1'b0;
    \A[588] = 1'b0;
    \A[589] = 1'b0;
    \A[590] = 1'b0;
    \A[591] = 1'b0;
    \A[592] = 1'b0;
    \A[593] = 1'b0;
    \A[594] = 1'b0;
    \A[595] = 1'b0;
    \A[596] = 1'b0;
    \A[597] = 1'b0;
    \A[598] = 1'b0;
    \A[599] = 1'b0;
    \A[600] = 1'b0;
    \A[601] = 1'b0;
    \A[602] = 1'b0;
    \A[603] = 1'b0;
    \A[604] = 1'b0;
    \A[605] = 1'b0;
    \A[606] = 1'b0;
    \A[607] = 1'b0;
    \A[608] = 1'b0;
    \A[609] = 1'b0;
    \A[610] = 1'b0;
    \A[611] = 1'b0;
    \A[612] = 1'b0;
    \A[613] = 1'b0;
    \A[614] = 1'b0;
    \A[615] = 1'b0;
    \A[616] = 1'b0;
    \A[617] = 1'b0;
    \A[618] = 1'b0;
    \A[619] = 1'b0;
    \A[620] = 1'b0;
    \A[621] = 1'b0;
    \A[622] = 1'b0;
    \A[623] = 1'b0;
    \A[624] = 1'b0;
    \A[625] = 1'b0;
    \A[626] = 1'b0;
    \A[627] = 1'b0;
    \A[628] = 1'b0;
    \A[629] = 1'b0;
    \A[630] = 1'b0;
    \A[631] = 1'b0;
    \A[632] = 1'b0;
    \A[633] = 1'b0;
    \A[634] = 1'b0;
    \A[635] = 1'b0;
    \A[636] = 1'b0;
    \A[637] = 1'b0;
    \A[638] = 1'b0;
    \A[639] = 1'b0;
    \A[640] = 1'b0;
    \A[641] = 1'b0;
    \A[642] = 1'b0;
    \A[643] = 1'b0;
    \A[644] = 1'b0;
    \A[645] = 1'b0;
    \A[646] = 1'b0;
    \A[647] = 1'b0;
    \A[648] = 1'b0;
    \A[649] = 1'b0;
    \A[650] = 1'b0;
    \A[651] = 1'b0;
    \A[652] = 1'b0;
    \A[653] = 1'b0;
    \A[654] = 1'b0;
    \A[655] = 1'b0;
    \A[656] = 1'b0;
    \A[657] = 1'b0;
    \A[658] = 1'b0;
    \A[659] = 1'b0;
    \A[660] = 1'b0;
    \A[661] = 1'b0;
    \A[662] = 1'b0;
    \A[663] = 1'b0;
    \A[664] = 1'b0;
    \A[665] = 1'b0;
    \A[666] = 1'b0;
    \A[667] = 1'b0;
    \A[668] = 1'b0;
    \A[669] = 1'b0;
    \A[670] = 1'b0;
    \A[671] = 1'b0;
    \A[672] = 1'b0;
    \A[673] = 1'b0;
    \A[674] = 1'b0;
    \A[675] = 1'b0;
    \A[676] = 1'b0;
    \A[677] = 1'b0;
    \A[678] = 1'b0;
    \A[679] = 1'b0;
    \A[680] = 1'b0;
    \A[681] = 1'b0;
    \A[682] = 1'b0;
    \A[683] = 1'b0;
    \A[684] = 1'b0;
    \A[685] = 1'b0;
    \A[686] = 1'b0;
    \A[687] = 1'b0;
    \A[688] = 1'b0;
    \A[689] = 1'b0;
    \A[690] = 1'b0;
    \A[691] = 1'b0;
    \A[692] = 1'b0;
    \A[693] = 1'b0;
    \A[694] = 1'b0;
    \A[695] = 1'b0;
    \A[696] = 1'b0;
    \A[697] = 1'b0;
    \A[698] = 1'b0;
    \A[699] = 1'b0;
    \A[700] = 1'b0;
    \A[701] = 1'b0;
    \A[702] = 1'b0;
    \A[703] = 1'b0;
    \A[704] = 1'b0;
    \A[705] = 1'b0;
    \A[706] = 1'b0;
    \A[707] = 1'b0;
    \A[708] = 1'b0;
    \A[709] = 1'b0;
    \A[710] = 1'b0;
    \A[711] = 1'b0;
    \A[712] = 1'b0;
    \A[713] = 1'b0;
    \A[714] = 1'b0;
    \A[715] = 1'b0;
    \A[716] = 1'b0;
    \A[717] = 1'b0;
    \A[718] = 1'b0;
    \A[719] = 1'b0;
    \A[720] = 1'b0;
    \A[721] = 1'b0;
    \A[722] = 1'b0;
    \A[723] = 1'b0;
    \A[724] = 1'b0;
    \A[725] = 1'b0;
    \A[726] = 1'b0;
    \A[727] = 1'b0;
    \A[728] = 1'b0;
    \A[729] = 1'b0;
    \A[730] = 1'b0;
    \A[731] = 1'b0;
    \A[732] = 1'b0;
    \A[733] = 1'b0;
    \A[734] = 1'b0;
    \A[735] = 1'b0;
    \A[736] = 1'b0;
    \A[737] = 1'b0;
    \A[738] = 1'b0;
    \A[739] = 1'b0;
    \A[740] = 1'b0;
    \A[741] = 1'b0;
    \A[742] = 1'b0;
    \A[743] = 1'b0;
    \A[744] = 1'b0;
    \A[745] = 1'b0;
    \A[746] = 1'b0;
    \A[747] = 1'b0;
    \A[748] = 1'b0;
    \A[749] = 1'b0;
    \A[750] = 1'b0;
    \A[751] = 1'b0;
    \A[752] = 1'b0;
    \A[753] = 1'b0;
    \A[754] = 1'b0;
    \A[755] = 1'b0;
    \A[756] = 1'b0;
    \A[757] = 1'b0;
    \A[758] = 1'b0;
    \A[759] = 1'b0;
    \A[760] = 1'b0;
    \A[761] = 1'b0;
    \A[762] = 1'b0;
    \A[763] = 1'b0;
    \A[764] = 1'b0;
    \A[765] = 1'b0;
    \A[766] = 1'b0;
    \A[767] = 1'b0;
    \A[768] = 1'b0;
    \A[769] = 1'b0;
    \A[770] = 1'b0;
    \A[771] = 1'b0;
    \A[772] = 1'b0;
    \A[773] = 1'b0;
    \A[774] = 1'b0;
    \A[775] = 1'b0;
    \A[776] = 1'b0;
    \A[777] = 1'b0;
    \A[778] = 1'b0;
    \A[779] = 1'b0;
    \A[780] = 1'b0;
    \A[781] = 1'b0;
    \A[782] = 1'b0;
    \A[783] = 1'b0;
    \A[784] = 1'b0;
    \A[785] = 1'b0;
    \A[786] = 1'b0;
    \A[787] = 1'b0;
    \A[788] = 1'b0;
    \A[789] = 1'b0;
    \A[790] = 1'b0;
    \A[791] = 1'b0;
    \A[792] = 1'b0;
    \A[793] = 1'b0;
    \A[794] = 1'b0;
    \A[795] = 1'b0;
    \A[796] = 1'b0;
    \A[797] = 1'b0;
    \A[798] = 1'b0;
    \A[799] = 1'b0;
    \A[800] = 1'b0;
    \A[801] = 1'b0;
    \A[802] = 1'b0;
    \A[803] = 1'b0;
    \A[804] = 1'b0;
    \A[805] = 1'b0;
    \A[806] = 1'b0;
    \A[807] = 1'b0;
    \A[808] = 1'b0;
    \A[809] = 1'b0;
    \A[810] = 1'b0;
    \A[811] = 1'b0;
    \A[812] = 1'b0;
    \A[813] = 1'b0;
    \A[814] = 1'b0;
    \A[815] = 1'b0;
    \A[816] = 1'b0;
    \A[817] = 1'b0;
    \A[818] = 1'b0;
    \A[819] = 1'b0;
    \A[820] = 1'b0;
    \A[821] = 1'b0;
    \A[822] = 1'b0;
    \A[823] = 1'b0;
    \A[824] = 1'b0;
    \A[825] = 1'b0;
    \A[826] = 1'b0;
    \A[827] = 1'b0;
    \A[828] = 1'b0;
    \A[829] = 1'b0;
    \A[830] = 1'b0;
    \A[831] = 1'b0;
    \A[832] = 1'b0;
    \A[833] = 1'b0;
    \A[834] = 1'b0;
    \A[835] = 1'b0;
    \A[836] = 1'b0;
    \A[837] = 1'b0;
    \A[838] = 1'b0;
    \A[839] = 1'b0;
    \A[840] = 1'b0;
    \A[841] = 1'b0;
    \A[842] = 1'b0;
    \A[843] = 1'b0;
    \A[844] = 1'b0;
    \A[845] = 1'b0;
    \A[846] = 1'b0;
    \A[847] = 1'b0;
    \A[848] = 1'b0;
    \A[849] = 1'b0;
    \A[850] = 1'b0;
    \A[851] = 1'b0;
    \A[852] = 1'b0;
    \A[853] = 1'b0;
    \A[854] = 1'b0;
    \A[855] = 1'b0;
    \A[856] = 1'b0;
    \A[857] = 1'b0;
    \A[858] = 1'b0;
    \A[859] = 1'b0;
    \A[860] = 1'b0;
    \A[861] = 1'b0;
    \A[862] = 1'b0;
    \A[863] = 1'b0;
    \A[864] = 1'b0;
    \A[865] = 1'b0;
    \A[866] = 1'b0;
    \A[867] = 1'b0;
    \A[868] = 1'b0;
    \A[869] = 1'b0;
    \A[870] = 1'b0;
    \A[871] = 1'b0;
    \A[872] = 1'b0;
    \A[873] = 1'b0;
    \A[874] = 1'b0;
    \A[875] = 1'b0;
    \A[876] = 1'b0;
    \A[877] = 1'b0;
    \A[878] = 1'b0;
    \A[879] = 1'b0;
    \A[880] = 1'b0;
    \A[881] = 1'b0;
    \A[882] = 1'b0;
    \A[883] = 1'b0;
    \A[884] = 1'b0;
    \A[885] = 1'b0;
    \A[886] = 1'b0;
    \A[887] = 1'b0;
    \A[888] = 1'b0;
    \A[889] = 1'b0;
    \A[890] = 1'b0;
    \A[891] = 1'b0;
    \A[892] = 1'b0;
    \A[893] = 1'b0;
    \A[894] = 1'b0;
    \A[895] = 1'b0;
    \A[896] = 1'b0;
    \A[897] = 1'b0;
    \A[898] = 1'b0;
    \A[899] = 1'b0;
    \A[900] = 1'b0;
    \A[901] = 1'b0;
    \A[902] = 1'b0;
    \A[903] = 1'b0;
    \A[904] = 1'b0;
    \A[905] = 1'b0;
    \A[906] = 1'b0;
    \A[907] = 1'b0;
    \A[908] = 1'b0;
    \A[909] = 1'b0;
    \A[910] = 1'b0;
    \A[911] = 1'b0;
    \A[912] = 1'b0;
    \A[913] = 1'b0;
    \A[914] = 1'b0;
    \A[915] = 1'b0;
    \A[916] = 1'b0;
    \A[917] = 1'b0;
    \A[918] = 1'b0;
    \A[919] = 1'b0;
    \A[920] = 1'b0;
    \A[921] = 1'b0;
    \A[922] = 1'b0;
    \A[923] = 1'b0;
    \A[924] = 1'b0;
    \A[925] = 1'b0;
    \A[926] = 1'b0;
    \A[927] = 1'b0;
    \A[928] = 1'b0;
    \A[929] = 1'b0;
    \A[930] = 1'b0;
    \A[931] = 1'b0;
    \A[932] = 1'b0;
    \A[933] = 1'b0;
    \A[934] = 1'b0;
    \A[935] = 1'b0;
    \A[936] = 1'b0;
    \A[937] = 1'b0;
    \A[938] = 1'b0;
    \A[939] = 1'b0;
    \A[940] = 1'b0;
    \A[941] = 1'b0;
    \A[942] = 1'b0;
    \A[943] = 1'b0;
    \A[944] = 1'b0;
    \A[945] = 1'b0;
    \A[946] = 1'b0;
    \A[947] = 1'b0;
    \A[948] = 1'b0;
    \A[949] = 1'b0;
    \A[950] = 1'b0;
    \A[951] = 1'b0;
    \A[952] = 1'b0;
    \A[953] = 1'b0;
    \A[954] = 1'b0;
    \A[955] = 1'b0;
    \A[956] = 1'b0;
    \A[957] = 1'b0;
    \A[958] = 1'b0;
    \A[959] = 1'b0;
    \A[960] = 1'b0;
    \A[961] = 1'b0;
    \A[962] = 1'b0;
    \A[963] = 1'b0;
    \A[964] = 1'b0;
    \A[965] = 1'b0;
    \A[966] = 1'b0;
    \A[967] = 1'b0;
    \A[968] = 1'b0;
    \A[969] = 1'b0;
    \A[970] = 1'b0;
    \A[971] = 1'b0;
    \A[972] = 1'b0;
    \A[973] = 1'b0;
    \A[974] = 1'b0;
    \A[975] = 1'b0;
    \A[976] = 1'b0;
    \A[977] = 1'b0;
    \A[978] = 1'b0;
    \A[979] = 1'b0;
    \A[980] = 1'b0;
    \A[981] = 1'b0;
    \A[982] = 1'b0;
    \A[983] = 1'b0;
    \A[984] = 1'b0;
    \A[985] = 1'b0;
    \A[986] = 1'b0;
    \A[987] = 1'b0;
    \A[988] = 1'b0;
    \A[989] = 1'b0;
    \A[990] = 1'b0;
    \A[991] = 1'b0;
    \A[992] = 1'b0;
    \A[993] = 1'b0;
    \A[994] = 1'b0;
    \A[995] = 1'b0;
    \A[996] = 1'b0;
    \A[997] = 1'b0;
    \A[998] = 1'b0;
    \A[999] = 1'b0;
    \A[1000] = 1'b0;

    #10;

    for (i = 0; i < STEPS; i = i + 1) begin

      // ===== 活跃区域激励 (64位) =====
      \A[0] = ((i / 2) % 2) ? 1'b1 : 1'b0;
      \A[1] = ((i / 4) % 2) ? 1'b1 : 1'b0;
      \A[2] = ((i / 8) % 2) ? 1'b1 : 1'b0;
      \A[3] = ((i / 16) % 2) ? 1'b1 : 1'b0;
      \A[4] = ((i / 32) % 2) ? 1'b1 : 1'b0;
      \A[5] = ((i / 64) % 2) ? 1'b1 : 1'b0;
      \A[6] = ((i / 128) % 2) ? 1'b1 : 1'b0;
      \A[7] = ((i / 256) % 2) ? 1'b1 : 1'b0;
      \A[8] = ((i / 2) % 2) ? 1'b1 : 1'b0;
      \A[9] = ((i / 4) % 2) ? 1'b1 : 1'b0;
      \A[10] = ((i / 8) % 2) ? 1'b1 : 1'b0;
      \A[11] = ((i / 16) % 2) ? 1'b1 : 1'b0;
      \A[12] = ((i / 32) % 2) ? 1'b1 : 1'b0;
      \A[13] = ((i / 64) % 2) ? 1'b1 : 1'b0;
      \A[14] = ((i / 128) % 2) ? 1'b1 : 1'b0;
      \A[15] = ((i / 256) % 2) ? 1'b1 : 1'b0;
      \A[16] = ((i / 2) % 2) ? 1'b1 : 1'b0;
      \A[17] = ((i / 4) % 2) ? 1'b1 : 1'b0;
      \A[18] = ((i / 8) % 2) ? 1'b1 : 1'b0;
      \A[19] = ((i / 16) % 2) ? 1'b1 : 1'b0;
      \A[20] = ((i / 32) % 2) ? 1'b1 : 1'b0;
      \A[21] = ((i / 64) % 2) ? 1'b1 : 1'b0;
      \A[22] = ((i / 128) % 2) ? 1'b1 : 1'b0;
      \A[23] = ((i / 256) % 2) ? 1'b1 : 1'b0;
      \A[24] = ((i / 2) % 2) ? 1'b1 : 1'b0;
      \A[25] = ((i / 4) % 2) ? 1'b1 : 1'b0;
      \A[26] = ((i / 8) % 2) ? 1'b1 : 1'b0;
      \A[27] = ((i / 16) % 2) ? 1'b1 : 1'b0;
      \A[28] = ((i / 32) % 2) ? 1'b1 : 1'b0;
      \A[29] = ((i / 64) % 2) ? 1'b1 : 1'b0;
      \A[30] = ((i / 128) % 2) ? 1'b1 : 1'b0;
      \A[31] = ((i / 256) % 2) ? 1'b1 : 1'b0;
      \A[32] = ((i / 2) % 2) ? 1'b1 : 1'b0;
      \A[33] = ((i / 4) % 2) ? 1'b1 : 1'b0;
      \A[34] = ((i / 8) % 2) ? 1'b1 : 1'b0;
      \A[35] = ((i / 16) % 2) ? 1'b1 : 1'b0;
      \A[36] = ((i / 32) % 2) ? 1'b1 : 1'b0;
      \A[37] = ((i / 64) % 2) ? 1'b1 : 1'b0;
      \A[38] = ((i / 128) % 2) ? 1'b1 : 1'b0;
      \A[39] = ((i / 256) % 2) ? 1'b1 : 1'b0;
      \A[40] = ((i / 2) % 2) ? 1'b1 : 1'b0;
      \A[41] = ((i / 4) % 2) ? 1'b1 : 1'b0;
      \A[42] = ((i / 8) % 2) ? 1'b1 : 1'b0;
      \A[43] = ((i / 16) % 2) ? 1'b1 : 1'b0;
      \A[44] = ((i / 32) % 2) ? 1'b1 : 1'b0;
      \A[45] = ((i / 64) % 2) ? 1'b1 : 1'b0;
      \A[46] = ((i / 128) % 2) ? 1'b1 : 1'b0;
      \A[47] = ((i / 256) % 2) ? 1'b1 : 1'b0;
      \A[48] = ((i / 2) % 2) ? 1'b1 : 1'b0;
      \A[49] = ((i / 4) % 2) ? 1'b1 : 1'b0;
      \A[50] = ((i / 8) % 2) ? 1'b1 : 1'b0;
      \A[51] = ((i / 16) % 2) ? 1'b1 : 1'b0;
      \A[52] = ((i / 32) % 2) ? 1'b1 : 1'b0;
      \A[53] = ((i / 64) % 2) ? 1'b1 : 1'b0;
      \A[54] = ((i / 128) % 2) ? 1'b1 : 1'b0;
      \A[55] = ((i / 256) % 2) ? 1'b1 : 1'b0;
      \A[56] = ((i / 2) % 2) ? 1'b1 : 1'b0;
      \A[57] = ((i / 4) % 2) ? 1'b1 : 1'b0;
      \A[58] = ((i / 8) % 2) ? 1'b1 : 1'b0;
      \A[59] = ((i / 16) % 2) ? 1'b1 : 1'b0;
      \A[60] = ((i / 32) % 2) ? 1'b1 : 1'b0;
      \A[61] = ((i / 64) % 2) ? 1'b1 : 1'b0;
      \A[62] = ((i / 128) % 2) ? 1'b1 : 1'b0;
      \A[63] = ((i / 256) % 2) ? 1'b1 : 1'b0;

      #10;

      if ((i % PRINT_EVERY) == 0) begin
        $display("o_sum=%06x", {maj});
      end
    end

    $display("o_sum=%06x [final]", {maj});
    $finish;
  end

  // VCD output
  reg [510:0] dumpfile_name;
  initial begin
    if (!$value$plusargs("DUMPFILE=%s", dumpfile_name)) begin
      $display("Error: No +DUMPFILE argument");
      $finish;
    end
    $display("Dumping VCD to: %s", dumpfile_name);
    $dumpfile(dumpfile_name);
    $dumpvars(0, tb);
  end

  initial begin
    #1;
    $display("FAULT_INJECTED: check_if_force_took_effect");
  end

endmodule