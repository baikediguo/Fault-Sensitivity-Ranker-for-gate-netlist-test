`timescale 1ns / 1ps

module tb;

  reg \A[0] ;
  reg \A[100] ;
  reg \A[101] ;
  reg \A[102] ;
  reg \A[103] ;
  reg \A[104] ;
  reg \A[105] ;
  reg \A[106] ;
  reg \A[107] ;
  reg \A[108] ;
  reg \A[109] ;
  reg \A[10] ;
  reg \A[110] ;
  reg \A[111] ;
  reg \A[112] ;
  reg \A[113] ;
  reg \A[114] ;
  reg \A[115] ;
  reg \A[116] ;
  reg \A[117] ;
  reg \A[118] ;
  reg \A[119] ;
  reg \A[11] ;
  reg \A[120] ;
  reg \A[121] ;
  reg \A[122] ;
  reg \A[123] ;
  reg \A[124] ;
  reg \A[125] ;
  reg \A[126] ;
  reg \A[127] ;
  reg \A[12] ;
  reg \A[13] ;
  reg \A[14] ;
  reg \A[15] ;
  reg \A[16] ;
  reg \A[17] ;
  reg \A[18] ;
  reg \A[19] ;
  reg \A[1] ;
  reg \A[20] ;
  reg \A[21] ;
  reg \A[22] ;
  reg \A[23] ;
  reg \A[24] ;
  reg \A[25] ;
  reg \A[26] ;
  reg \A[27] ;
  reg \A[28] ;
  reg \A[29] ;
  reg \A[2] ;
  reg \A[30] ;
  reg \A[31] ;
  reg \A[32] ;
  reg \A[33] ;
  reg \A[34] ;
  reg \A[35] ;
  reg \A[36] ;
  reg \A[37] ;
  reg \A[38] ;
  reg \A[39] ;
  reg \A[3] ;
  reg \A[40] ;
  reg \A[41] ;
  reg \A[42] ;
  reg \A[43] ;
  reg \A[44] ;
  reg \A[45] ;
  reg \A[46] ;
  reg \A[47] ;
  reg \A[48] ;
  reg \A[49] ;
  reg \A[4] ;
  reg \A[50] ;
  reg \A[51] ;
  reg \A[52] ;
  reg \A[53] ;
  reg \A[54] ;
  reg \A[55] ;
  reg \A[56] ;
  reg \A[57] ;
  reg \A[58] ;
  reg \A[59] ;
  reg \A[5] ;
  reg \A[60] ;
  reg \A[61] ;
  reg \A[62] ;
  reg \A[63] ;
  reg \A[64] ;
  reg \A[65] ;
  reg \A[66] ;
  reg \A[67] ;
  reg \A[68] ;
  reg \A[69] ;
  reg \A[6] ;
  reg \A[70] ;
  reg \A[71] ;
  reg \A[72] ;
  reg \A[73] ;
  reg \A[74] ;
  reg \A[75] ;
  reg \A[76] ;
  reg \A[77] ;
  reg \A[78] ;
  reg \A[79] ;
  reg \A[7] ;
  reg \A[80] ;
  reg \A[81] ;
  reg \A[82] ;
  reg \A[83] ;
  reg \A[84] ;
  reg \A[85] ;
  reg \A[86] ;
  reg \A[87] ;
  reg \A[88] ;
  reg \A[89] ;
  reg \A[8] ;
  reg \A[90] ;
  reg \A[91] ;
  reg \A[92] ;
  reg \A[93] ;
  reg \A[94] ;
  reg \A[95] ;
  reg \A[96] ;
  reg \A[97] ;
  reg \A[98] ;
  reg \A[99] ;
  reg \A[9] ;
  wire \P[0] ;
  wire \P[1] ;
  wire \P[2] ;
  wire \P[3] ;
  wire \P[4] ;
  wire \P[5] ;
  wire \P[6] ;
  wire F;

  // DUT (combinational)
  top uut (
    .\A[0] (\A[0] ),
    .\A[100] (\A[100] ),
    .\A[101] (\A[101] ),
    .\A[102] (\A[102] ),
    .\A[103] (\A[103] ),
    .\A[104] (\A[104] ),
    .\A[105] (\A[105] ),
    .\A[106] (\A[106] ),
    .\A[107] (\A[107] ),
    .\A[108] (\A[108] ),
    .\A[109] (\A[109] ),
    .\A[10] (\A[10] ),
    .\A[110] (\A[110] ),
    .\A[111] (\A[111] ),
    .\A[112] (\A[112] ),
    .\A[113] (\A[113] ),
    .\A[114] (\A[114] ),
    .\A[115] (\A[115] ),
    .\A[116] (\A[116] ),
    .\A[117] (\A[117] ),
    .\A[118] (\A[118] ),
    .\A[119] (\A[119] ),
    .\A[11] (\A[11] ),
    .\A[120] (\A[120] ),
    .\A[121] (\A[121] ),
    .\A[122] (\A[122] ),
    .\A[123] (\A[123] ),
    .\A[124] (\A[124] ),
    .\A[125] (\A[125] ),
    .\A[126] (\A[126] ),
    .\A[127] (\A[127] ),
    .\A[12] (\A[12] ),
    .\A[13] (\A[13] ),
    .\A[14] (\A[14] ),
    .\A[15] (\A[15] ),
    .\A[16] (\A[16] ),
    .\A[17] (\A[17] ),
    .\A[18] (\A[18] ),
    .\A[19] (\A[19] ),
    .\A[1] (\A[1] ),
    .\A[20] (\A[20] ),
    .\A[21] (\A[21] ),
    .\A[22] (\A[22] ),
    .\A[23] (\A[23] ),
    .\A[24] (\A[24] ),
    .\A[25] (\A[25] ),
    .\A[26] (\A[26] ),
    .\A[27] (\A[27] ),
    .\A[28] (\A[28] ),
    .\A[29] (\A[29] ),
    .\A[2] (\A[2] ),
    .\A[30] (\A[30] ),
    .\A[31] (\A[31] ),
    .\A[32] (\A[32] ),
    .\A[33] (\A[33] ),
    .\A[34] (\A[34] ),
    .\A[35] (\A[35] ),
    .\A[36] (\A[36] ),
    .\A[37] (\A[37] ),
    .\A[38] (\A[38] ),
    .\A[39] (\A[39] ),
    .\A[3] (\A[3] ),
    .\A[40] (\A[40] ),
    .\A[41] (\A[41] ),
    .\A[42] (\A[42] ),
    .\A[43] (\A[43] ),
    .\A[44] (\A[44] ),
    .\A[45] (\A[45] ),
    .\A[46] (\A[46] ),
    .\A[47] (\A[47] ),
    .\A[48] (\A[48] ),
    .\A[49] (\A[49] ),
    .\A[4] (\A[4] ),
    .\A[50] (\A[50] ),
    .\A[51] (\A[51] ),
    .\A[52] (\A[52] ),
    .\A[53] (\A[53] ),
    .\A[54] (\A[54] ),
    .\A[55] (\A[55] ),
    .\A[56] (\A[56] ),
    .\A[57] (\A[57] ),
    .\A[58] (\A[58] ),
    .\A[59] (\A[59] ),
    .\A[5] (\A[5] ),
    .\A[60] (\A[60] ),
    .\A[61] (\A[61] ),
    .\A[62] (\A[62] ),
    .\A[63] (\A[63] ),
    .\A[64] (\A[64] ),
    .\A[65] (\A[65] ),
    .\A[66] (\A[66] ),
    .\A[67] (\A[67] ),
    .\A[68] (\A[68] ),
    .\A[69] (\A[69] ),
    .\A[6] (\A[6] ),
    .\A[70] (\A[70] ),
    .\A[71] (\A[71] ),
    .\A[72] (\A[72] ),
    .\A[73] (\A[73] ),
    .\A[74] (\A[74] ),
    .\A[75] (\A[75] ),
    .\A[76] (\A[76] ),
    .\A[77] (\A[77] ),
    .\A[78] (\A[78] ),
    .\A[79] (\A[79] ),
    .\A[7] (\A[7] ),
    .\A[80] (\A[80] ),
    .\A[81] (\A[81] ),
    .\A[82] (\A[82] ),
    .\A[83] (\A[83] ),
    .\A[84] (\A[84] ),
    .\A[85] (\A[85] ),
    .\A[86] (\A[86] ),
    .\A[87] (\A[87] ),
    .\A[88] (\A[88] ),
    .\A[89] (\A[89] ),
    .\A[8] (\A[8] ),
    .\A[90] (\A[90] ),
    .\A[91] (\A[91] ),
    .\A[92] (\A[92] ),
    .\A[93] (\A[93] ),
    .\A[94] (\A[94] ),
    .\A[95] (\A[95] ),
    .\A[96] (\A[96] ),
    .\A[97] (\A[97] ),
    .\A[98] (\A[98] ),
    .\A[99] (\A[99] ),
    .\A[9] (\A[9] ),
    .\P[0] (\P[0] ),
    .\P[1] (\P[1] ),
    .\P[2] (\P[2] ),
    .\P[3] (\P[3] ),
    .\P[4] (\P[4] ),
    .\P[5] (\P[5] ),
    .\P[6] (\P[6] ),
    .F(F)
  );

  // Random function
  integer SEED = 6;
  function [7:0] urand(input integer s);
    urand = $random(s) & 8'hFF;
  endfunction

  // Main stimulus (combinational)
  integer i;
  parameter CYCLES = 512;
  parameter PRINT_EVERY = 1;

  initial begin
    \A[0] = 0;
    \A[100] = 0;
    \A[101] = 0;
    \A[102] = 0;
    \A[103] = 0;
    \A[104] = 0;
    \A[105] = 0;
    \A[106] = 0;
    \A[107] = 0;
    \A[108] = 0;
    \A[109] = 0;
    \A[10] = 0;
    \A[110] = 0;
    \A[111] = 0;
    \A[112] = 0;
    \A[113] = 0;
    \A[114] = 0;
    \A[115] = 0;
    \A[116] = 0;
    \A[117] = 0;
    \A[118] = 0;
    \A[119] = 0;
    \A[11] = 0;
    \A[120] = 0;
    \A[121] = 0;
    \A[122] = 0;
    \A[123] = 0;
    \A[124] = 0;
    \A[125] = 0;
    \A[126] = 0;
    \A[127] = 0;
    \A[12] = 0;
    \A[13] = 0;
    \A[14] = 0;
    \A[15] = 0;
    \A[16] = 0;
    \A[17] = 0;
    \A[18] = 0;
    \A[19] = 0;
    \A[1] = 0;
    \A[20] = 0;
    \A[21] = 0;
    \A[22] = 0;
    \A[23] = 0;
    \A[24] = 0;
    \A[25] = 0;
    \A[26] = 0;
    \A[27] = 0;
    \A[28] = 0;
    \A[29] = 0;
    \A[2] = 0;
    \A[30] = 0;
    \A[31] = 0;
    \A[32] = 0;
    \A[33] = 0;
    \A[34] = 0;
    \A[35] = 0;
    \A[36] = 0;
    \A[37] = 0;
    \A[38] = 0;
    \A[39] = 0;
    \A[3] = 0;
    \A[40] = 0;
    \A[41] = 0;
    \A[42] = 0;
    \A[43] = 0;
    \A[44] = 0;
    \A[45] = 0;
    \A[46] = 0;
    \A[47] = 0;
    \A[48] = 0;
    \A[49] = 0;
    \A[4] = 0;
    \A[50] = 0;
    \A[51] = 0;
    \A[52] = 0;
    \A[53] = 0;
    \A[54] = 0;
    \A[55] = 0;
    \A[56] = 0;
    \A[57] = 0;
    \A[58] = 0;
    \A[59] = 0;
    \A[5] = 0;
    \A[60] = 0;
    \A[61] = 0;
    \A[62] = 0;
    \A[63] = 0;
    \A[64] = 0;
    \A[65] = 0;
    \A[66] = 0;
    \A[67] = 0;
    \A[68] = 0;
    \A[69] = 0;
    \A[6] = 0;
    \A[70] = 0;
    \A[71] = 0;
    \A[72] = 0;
    \A[73] = 0;
    \A[74] = 0;
    \A[75] = 0;
    \A[76] = 0;
    \A[77] = 0;
    \A[78] = 0;
    \A[79] = 0;
    \A[7] = 0;
    \A[80] = 0;
    \A[81] = 0;
    \A[82] = 0;
    \A[83] = 0;
    \A[84] = 0;
    \A[85] = 0;
    \A[86] = 0;
    \A[87] = 0;
    \A[88] = 0;
    \A[89] = 0;
    \A[8] = 0;
    \A[90] = 0;
    \A[91] = 0;
    \A[92] = 0;
    \A[93] = 0;
    \A[94] = 0;
    \A[95] = 0;
    \A[96] = 0;
    \A[97] = 0;
    \A[98] = 0;
    \A[99] = 0;
    \A[9] = 0;

    #10;

    for (i = 0; i < CYCLES; i = i + 1) begin
        // \A[0]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[0] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[0] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[0] = (i + 0) % 2;  // Phase3: 翻转
          end
        end

        // \A[100]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[100] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[100] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[100] = (i + 1) % 2;  // Phase3: 翻转
          end
        end

        // \A[101]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[101] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[101] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[101] = (i + 2) % 2;  // Phase3: 翻转
          end
        end

        // \A[102]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[102] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[102] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[102] = (i + 3) % 2;  // Phase3: 翻转
          end
        end

        // \A[103]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[103] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[103] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[103] = (i + 4) % 2;  // Phase3: 翻转
          end
        end

        // \A[104]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[104] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[104] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[104] = (i + 5) % 2;  // Phase3: 翻转
          end
        end

        // \A[105]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[105] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[105] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[105] = (i + 6) % 2;  // Phase3: 翻转
          end
        end

        // \A[106]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[106] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[106] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[106] = (i + 7) % 2;  // Phase3: 翻转
          end
        end

        // \A[107]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[107] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[107] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[107] = (i + 8) % 2;  // Phase3: 翻转
          end
        end

        // \A[108]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[108] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[108] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[108] = (i + 9) % 2;  // Phase3: 翻转
          end
        end

        // \A[109]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[109] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[109] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[109] = (i + 10) % 2;  // Phase3: 翻转
          end
        end

        // \A[10]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[10] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[10] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[10] = (i + 11) % 2;  // Phase3: 翻转
          end
        end

        // \A[110]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[110] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[110] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[110] = (i + 12) % 2;  // Phase3: 翻转
          end
        end

        // \A[111]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[111] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[111] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[111] = (i + 13) % 2;  // Phase3: 翻转
          end
        end

        // \A[112]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[112] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[112] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[112] = (i + 14) % 2;  // Phase3: 翻转
          end
        end

        // \A[113]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[113] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[113] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[113] = (i + 15) % 2;  // Phase3: 翻转
          end
        end

        // \A[114]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[114] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[114] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[114] = (i + 16) % 2;  // Phase3: 翻转
          end
        end

        // \A[115]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[115] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[115] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[115] = (i + 17) % 2;  // Phase3: 翻转
          end
        end

        // \A[116]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[116] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[116] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[116] = (i + 18) % 2;  // Phase3: 翻转
          end
        end

        // \A[117]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[117] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[117] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[117] = (i + 19) % 2;  // Phase3: 翻转
          end
        end

        // \A[118]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[118] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[118] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[118] = (i + 20) % 2;  // Phase3: 翻转
          end
        end

        // \A[119]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[119] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[119] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[119] = (i + 21) % 2;  // Phase3: 翻转
          end
        end

        // \A[11]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[11] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[11] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[11] = (i + 22) % 2;  // Phase3: 翻转
          end
        end

        // \A[120]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[120] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[120] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[120] = (i + 23) % 2;  // Phase3: 翻转
          end
        end

        // \A[121]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[121] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[121] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[121] = (i + 24) % 2;  // Phase3: 翻转
          end
        end

        // \A[122]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[122] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[122] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[122] = (i + 25) % 2;  // Phase3: 翻转
          end
        end

        // \A[123]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[123] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[123] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[123] = (i + 26) % 2;  // Phase3: 翻转
          end
        end

        // \A[124]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[124] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[124] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[124] = (i + 27) % 2;  // Phase3: 翻转
          end
        end

        // \A[125]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[125] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[125] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[125] = (i + 28) % 2;  // Phase3: 翻转
          end
        end

        // \A[126]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[126] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[126] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[126] = (i + 29) % 2;  // Phase3: 翻转
          end
        end

        // \A[127]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[127] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[127] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[127] = (i + 30) % 2;  // Phase3: 翻转
          end
        end

        // \A[12]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[12] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[12] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[12] = (i + 31) % 2;  // Phase3: 翻转
          end
        end

        // \A[13]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[13] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[13] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[13] = (i + 32) % 2;  // Phase3: 翻转
          end
        end

        // \A[14]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[14] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[14] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[14] = (i + 33) % 2;  // Phase3: 翻转
          end
        end

        // \A[15]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[15] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[15] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[15] = (i + 34) % 2;  // Phase3: 翻转
          end
        end

        // \A[16]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[16] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[16] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[16] = (i + 35) % 2;  // Phase3: 翻转
          end
        end

        // \A[17]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[17] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[17] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[17] = (i + 36) % 2;  // Phase3: 翻转
          end
        end

        // \A[18]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[18] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[18] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[18] = (i + 37) % 2;  // Phase3: 翻转
          end
        end

        // \A[19]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[19] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[19] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[19] = (i + 38) % 2;  // Phase3: 翻转
          end
        end

        // \A[1]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[1] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[1] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[1] = (i + 39) % 2;  // Phase3: 翻转
          end
        end

        // \A[20]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[20] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[20] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[20] = (i + 40) % 2;  // Phase3: 翻转
          end
        end

        // \A[21]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[21] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[21] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[21] = (i + 41) % 2;  // Phase3: 翻转
          end
        end

        // \A[22]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[22] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[22] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[22] = (i + 42) % 2;  // Phase3: 翻转
          end
        end

        // \A[23]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[23] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[23] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[23] = (i + 43) % 2;  // Phase3: 翻转
          end
        end

        // \A[24]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[24] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[24] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[24] = (i + 44) % 2;  // Phase3: 翻转
          end
        end

        // \A[25]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[25] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[25] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[25] = (i + 45) % 2;  // Phase3: 翻转
          end
        end

        // \A[26]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[26] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[26] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[26] = (i + 46) % 2;  // Phase3: 翻转
          end
        end

        // \A[27]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[27] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[27] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[27] = (i + 47) % 2;  // Phase3: 翻转
          end
        end

        // \A[28]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[28] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[28] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[28] = (i + 48) % 2;  // Phase3: 翻转
          end
        end

        // \A[29]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[29] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[29] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[29] = (i + 49) % 2;  // Phase3: 翻转
          end
        end

        // \A[2]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[2] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[2] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[2] = (i + 50) % 2;  // Phase3: 翻转
          end
        end

        // \A[30]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[30] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[30] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[30] = (i + 51) % 2;  // Phase3: 翻转
          end
        end

        // \A[31]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[31] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[31] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[31] = (i + 52) % 2;  // Phase3: 翻转
          end
        end

        // \A[32]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[32] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[32] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[32] = (i + 53) % 2;  // Phase3: 翻转
          end
        end

        // \A[33]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[33] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[33] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[33] = (i + 54) % 2;  // Phase3: 翻转
          end
        end

        // \A[34]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[34] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[34] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[34] = (i + 55) % 2;  // Phase3: 翻转
          end
        end

        // \A[35]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[35] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[35] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[35] = (i + 56) % 2;  // Phase3: 翻转
          end
        end

        // \A[36]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[36] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[36] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[36] = (i + 57) % 2;  // Phase3: 翻转
          end
        end

        // \A[37]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[37] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[37] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[37] = (i + 58) % 2;  // Phase3: 翻转
          end
        end

        // \A[38]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[38] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[38] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[38] = (i + 59) % 2;  // Phase3: 翻转
          end
        end

        // \A[39]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[39] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[39] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[39] = (i + 60) % 2;  // Phase3: 翻转
          end
        end

        // \A[3]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[3] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[3] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[3] = (i + 61) % 2;  // Phase3: 翻转
          end
        end

        // \A[40]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[40] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[40] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[40] = (i + 62) % 2;  // Phase3: 翻转
          end
        end

        // \A[41]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[41] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[41] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[41] = (i + 63) % 2;  // Phase3: 翻转
          end
        end

        // \A[42]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[42] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[42] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[42] = (i + 64) % 2;  // Phase3: 翻转
          end
        end

        // \A[43]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[43] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[43] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[43] = (i + 65) % 2;  // Phase3: 翻转
          end
        end

        // \A[44]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[44] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[44] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[44] = (i + 66) % 2;  // Phase3: 翻转
          end
        end

        // \A[45]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[45] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[45] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[45] = (i + 67) % 2;  // Phase3: 翻转
          end
        end

        // \A[46]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[46] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[46] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[46] = (i + 68) % 2;  // Phase3: 翻转
          end
        end

        // \A[47]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[47] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[47] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[47] = (i + 69) % 2;  // Phase3: 翻转
          end
        end

        // \A[48]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[48] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[48] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[48] = (i + 70) % 2;  // Phase3: 翻转
          end
        end

        // \A[49]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[49] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[49] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[49] = (i + 71) % 2;  // Phase3: 翻转
          end
        end

        // \A[4]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[4] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[4] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[4] = (i + 72) % 2;  // Phase3: 翻转
          end
        end

        // \A[50]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[50] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[50] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[50] = (i + 73) % 2;  // Phase3: 翻转
          end
        end

        // \A[51]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[51] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[51] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[51] = (i + 74) % 2;  // Phase3: 翻转
          end
        end

        // \A[52]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[52] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[52] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[52] = (i + 75) % 2;  // Phase3: 翻转
          end
        end

        // \A[53]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[53] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[53] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[53] = (i + 76) % 2;  // Phase3: 翻转
          end
        end

        // \A[54]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[54] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[54] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[54] = (i + 77) % 2;  // Phase3: 翻转
          end
        end

        // \A[55]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[55] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[55] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[55] = (i + 78) % 2;  // Phase3: 翻转
          end
        end

        // \A[56]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[56] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[56] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[56] = (i + 79) % 2;  // Phase3: 翻转
          end
        end

        // \A[57]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[57] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[57] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[57] = (i + 80) % 2;  // Phase3: 翻转
          end
        end

        // \A[58]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[58] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[58] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[58] = (i + 81) % 2;  // Phase3: 翻转
          end
        end

        // \A[59]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[59] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[59] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[59] = (i + 82) % 2;  // Phase3: 翻转
          end
        end

        // \A[5]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[5] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[5] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[5] = (i + 83) % 2;  // Phase3: 翻转
          end
        end

        // \A[60]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[60] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[60] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[60] = (i + 84) % 2;  // Phase3: 翻转
          end
        end

        // \A[61]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[61] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[61] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[61] = (i + 85) % 2;  // Phase3: 翻转
          end
        end

        // \A[62]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[62] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[62] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[62] = (i + 86) % 2;  // Phase3: 翻转
          end
        end

        // \A[63]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[63] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[63] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[63] = (i + 87) % 2;  // Phase3: 翻转
          end
        end

        // \A[64]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[64] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[64] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[64] = (i + 88) % 2;  // Phase3: 翻转
          end
        end

        // \A[65]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[65] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[65] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[65] = (i + 89) % 2;  // Phase3: 翻转
          end
        end

        // \A[66]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[66] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[66] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[66] = (i + 90) % 2;  // Phase3: 翻转
          end
        end

        // \A[67]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[67] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[67] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[67] = (i + 91) % 2;  // Phase3: 翻转
          end
        end

        // \A[68]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[68] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[68] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[68] = (i + 92) % 2;  // Phase3: 翻转
          end
        end

        // \A[69]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[69] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[69] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[69] = (i + 93) % 2;  // Phase3: 翻转
          end
        end

        // \A[6]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[6] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[6] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[6] = (i + 94) % 2;  // Phase3: 翻转
          end
        end

        // \A[70]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[70] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[70] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[70] = (i + 95) % 2;  // Phase3: 翻转
          end
        end

        // \A[71]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[71] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[71] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[71] = (i + 96) % 2;  // Phase3: 翻转
          end
        end

        // \A[72]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[72] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[72] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[72] = (i + 97) % 2;  // Phase3: 翻转
          end
        end

        // \A[73]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[73] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[73] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[73] = (i + 98) % 2;  // Phase3: 翻转
          end
        end

        // \A[74]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[74] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[74] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[74] = (i + 99) % 2;  // Phase3: 翻转
          end
        end

        // \A[75]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[75] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[75] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[75] = (i + 100) % 2;  // Phase3: 翻转
          end
        end

        // \A[76]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[76] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[76] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[76] = (i + 101) % 2;  // Phase3: 翻转
          end
        end

        // \A[77]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[77] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[77] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[77] = (i + 102) % 2;  // Phase3: 翻转
          end
        end

        // \A[78]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[78] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[78] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[78] = (i + 103) % 2;  // Phase3: 翻转
          end
        end

        // \A[79]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[79] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[79] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[79] = (i + 104) % 2;  // Phase3: 翻转
          end
        end

        // \A[7]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[7] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[7] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[7] = (i + 105) % 2;  // Phase3: 翻转
          end
        end

        // \A[80]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[80] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[80] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[80] = (i + 106) % 2;  // Phase3: 翻转
          end
        end

        // \A[81]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[81] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[81] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[81] = (i + 107) % 2;  // Phase3: 翻转
          end
        end

        // \A[82]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[82] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[82] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[82] = (i + 108) % 2;  // Phase3: 翻转
          end
        end

        // \A[83]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[83] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[83] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[83] = (i + 109) % 2;  // Phase3: 翻转
          end
        end

        // \A[84]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[84] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[84] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[84] = (i + 110) % 2;  // Phase3: 翻转
          end
        end

        // \A[85]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[85] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[85] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[85] = (i + 111) % 2;  // Phase3: 翻转
          end
        end

        // \A[86]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[86] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[86] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[86] = (i + 112) % 2;  // Phase3: 翻转
          end
        end

        // \A[87]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[87] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[87] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[87] = (i + 113) % 2;  // Phase3: 翻转
          end
        end

        // \A[88]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[88] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[88] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[88] = (i + 114) % 2;  // Phase3: 翻转
          end
        end

        // \A[89]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[89] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[89] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[89] = (i + 115) % 2;  // Phase3: 翻转
          end
        end

        // \A[8]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[8] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[8] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[8] = (i + 116) % 2;  // Phase3: 翻转
          end
        end

        // \A[90]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[90] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[90] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[90] = (i + 117) % 2;  // Phase3: 翻转
          end
        end

        // \A[91]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[91] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[91] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[91] = (i + 118) % 2;  // Phase3: 翻转
          end
        end

        // \A[92]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[92] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[92] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[92] = (i + 119) % 2;  // Phase3: 翻转
          end
        end

        // \A[93]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[93] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[93] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[93] = (i + 120) % 2;  // Phase3: 翻转
          end
        end

        // \A[94]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[94] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[94] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[94] = (i + 121) % 2;  // Phase3: 翻转
          end
        end

        // \A[95]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[95] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[95] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[95] = (i + 122) % 2;  // Phase3: 翻转
          end
        end

        // \A[96]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[96] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[96] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[96] = (i + 123) % 2;  // Phase3: 翻转
          end
        end

        // \A[97]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[97] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[97] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[97] = (i + 124) % 2;  // Phase3: 翻转
          end
        end

        // \A[98]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[98] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[98] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[98] = (i + 125) % 2;  // Phase3: 翻转
          end
        end

        // \A[99]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[99] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[99] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[99] = (i + 126) % 2;  // Phase3: 翻转
          end
        end

        // \A[9]: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            \A[9] = 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            \A[9] = 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            \A[9] = (i + 127) % 2;  // Phase3: 翻转
          end
        end

      #10;

      if ((i % PRINT_EVERY) == 0) begin
        $display("o_sum=%06x", {\P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F});
      end
    end

    $display("o_sum=%06x [final]", {\P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F});
    $finish;
  end

  // VCD output (optional)
  reg [510:0] dumpfile_name;
  initial begin
    if ($value$plusargs("DUMPFILE=%s", dumpfile_name)) begin
      $display("Dumping VCD to: %s", dumpfile_name);
      $dumpfile(dumpfile_name);
      $dumpvars(0, tb);
    end
  end

  initial begin
    #1;
    $display("FAULT_INJECTED: check_if_force_took_effect");
  end

endmodule
