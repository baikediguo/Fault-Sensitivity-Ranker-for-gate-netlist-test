`timescale 1ns / 1ps

module tb;

  reg [127:0] a_vec;
  reg [127:0] b_vec;
  wire [127:0] hyp_vec;

  top uut (
    .\a[0] (a_vec[0]),     .\a[1] (a_vec[1]),     .\a[2] (a_vec[2]),     .\a[3] (a_vec[3]),     .\a[4] (a_vec[4]),     .\a[5] (a_vec[5]),     .\a[6] (a_vec[6]),     .\a[7] (a_vec[7]), 
    .\a[8] (a_vec[8]),     .\a[9] (a_vec[9]),     .\a[10] (a_vec[10]),     .\a[11] (a_vec[11]),     .\a[12] (a_vec[12]),     .\a[13] (a_vec[13]),     .\a[14] (a_vec[14]),     .\a[15] (a_vec[15]), 
    .\a[16] (a_vec[16]),     .\a[17] (a_vec[17]),     .\a[18] (a_vec[18]),     .\a[19] (a_vec[19]),     .\a[20] (a_vec[20]),     .\a[21] (a_vec[21]),     .\a[22] (a_vec[22]),     .\a[23] (a_vec[23]), 
    .\a[24] (a_vec[24]),     .\a[25] (a_vec[25]),     .\a[26] (a_vec[26]),     .\a[27] (a_vec[27]),     .\a[28] (a_vec[28]),     .\a[29] (a_vec[29]),     .\a[30] (a_vec[30]),     .\a[31] (a_vec[31]), 
    .\a[32] (a_vec[32]),     .\a[33] (a_vec[33]),     .\a[34] (a_vec[34]),     .\a[35] (a_vec[35]),     .\a[36] (a_vec[36]),     .\a[37] (a_vec[37]),     .\a[38] (a_vec[38]),     .\a[39] (a_vec[39]), 
    .\a[40] (a_vec[40]),     .\a[41] (a_vec[41]),     .\a[42] (a_vec[42]),     .\a[43] (a_vec[43]),     .\a[44] (a_vec[44]),     .\a[45] (a_vec[45]),     .\a[46] (a_vec[46]),     .\a[47] (a_vec[47]), 
    .\a[48] (a_vec[48]),     .\a[49] (a_vec[49]),     .\a[50] (a_vec[50]),     .\a[51] (a_vec[51]),     .\a[52] (a_vec[52]),     .\a[53] (a_vec[53]),     .\a[54] (a_vec[54]),     .\a[55] (a_vec[55]), 
    .\a[56] (a_vec[56]),     .\a[57] (a_vec[57]),     .\a[58] (a_vec[58]),     .\a[59] (a_vec[59]),     .\a[60] (a_vec[60]),     .\a[61] (a_vec[61]),     .\a[62] (a_vec[62]),     .\a[63] (a_vec[63]), 
    .\a[64] (a_vec[64]),     .\a[65] (a_vec[65]),     .\a[66] (a_vec[66]),     .\a[67] (a_vec[67]),     .\a[68] (a_vec[68]),     .\a[69] (a_vec[69]),     .\a[70] (a_vec[70]),     .\a[71] (a_vec[71]), 
    .\a[72] (a_vec[72]),     .\a[73] (a_vec[73]),     .\a[74] (a_vec[74]),     .\a[75] (a_vec[75]),     .\a[76] (a_vec[76]),     .\a[77] (a_vec[77]),     .\a[78] (a_vec[78]),     .\a[79] (a_vec[79]), 
    .\a[80] (a_vec[80]),     .\a[81] (a_vec[81]),     .\a[82] (a_vec[82]),     .\a[83] (a_vec[83]),     .\a[84] (a_vec[84]),     .\a[85] (a_vec[85]),     .\a[86] (a_vec[86]),     .\a[87] (a_vec[87]), 
    .\a[88] (a_vec[88]),     .\a[89] (a_vec[89]),     .\a[90] (a_vec[90]),     .\a[91] (a_vec[91]),     .\a[92] (a_vec[92]),     .\a[93] (a_vec[93]),     .\a[94] (a_vec[94]),     .\a[95] (a_vec[95]), 
    .\a[96] (a_vec[96]),     .\a[97] (a_vec[97]),     .\a[98] (a_vec[98]),     .\a[99] (a_vec[99]),     .\a[100] (a_vec[100]),     .\a[101] (a_vec[101]),     .\a[102] (a_vec[102]),     .\a[103] (a_vec[103]), 
    .\a[104] (a_vec[104]),     .\a[105] (a_vec[105]),     .\a[106] (a_vec[106]),     .\a[107] (a_vec[107]),     .\a[108] (a_vec[108]),     .\a[109] (a_vec[109]),     .\a[110] (a_vec[110]),     .\a[111] (a_vec[111]), 
    .\a[112] (a_vec[112]),     .\a[113] (a_vec[113]),     .\a[114] (a_vec[114]),     .\a[115] (a_vec[115]),     .\a[116] (a_vec[116]),     .\a[117] (a_vec[117]),     .\a[118] (a_vec[118]),     .\a[119] (a_vec[119]), 
    .\a[120] (a_vec[120]),     .\a[121] (a_vec[121]),     .\a[122] (a_vec[122]),     .\a[123] (a_vec[123]),     .\a[124] (a_vec[124]),     .\a[125] (a_vec[125]),     .\a[126] (a_vec[126]),     .\a[127] (a_vec[127]), 
    .\b[0] (b_vec[0]),     .\b[1] (b_vec[1]),     .\b[2] (b_vec[2]),     .\b[3] (b_vec[3]),     .\b[4] (b_vec[4]),     .\b[5] (b_vec[5]),     .\b[6] (b_vec[6]),     .\b[7] (b_vec[7]), 
    .\b[8] (b_vec[8]),     .\b[9] (b_vec[9]),     .\b[10] (b_vec[10]),     .\b[11] (b_vec[11]),     .\b[12] (b_vec[12]),     .\b[13] (b_vec[13]),     .\b[14] (b_vec[14]),     .\b[15] (b_vec[15]), 
    .\b[16] (b_vec[16]),     .\b[17] (b_vec[17]),     .\b[18] (b_vec[18]),     .\b[19] (b_vec[19]),     .\b[20] (b_vec[20]),     .\b[21] (b_vec[21]),     .\b[22] (b_vec[22]),     .\b[23] (b_vec[23]), 
    .\b[24] (b_vec[24]),     .\b[25] (b_vec[25]),     .\b[26] (b_vec[26]),     .\b[27] (b_vec[27]),     .\b[28] (b_vec[28]),     .\b[29] (b_vec[29]),     .\b[30] (b_vec[30]),     .\b[31] (b_vec[31]), 
    .\b[32] (b_vec[32]),     .\b[33] (b_vec[33]),     .\b[34] (b_vec[34]),     .\b[35] (b_vec[35]),     .\b[36] (b_vec[36]),     .\b[37] (b_vec[37]),     .\b[38] (b_vec[38]),     .\b[39] (b_vec[39]), 
    .\b[40] (b_vec[40]),     .\b[41] (b_vec[41]),     .\b[42] (b_vec[42]),     .\b[43] (b_vec[43]),     .\b[44] (b_vec[44]),     .\b[45] (b_vec[45]),     .\b[46] (b_vec[46]),     .\b[47] (b_vec[47]), 
    .\b[48] (b_vec[48]),     .\b[49] (b_vec[49]),     .\b[50] (b_vec[50]),     .\b[51] (b_vec[51]),     .\b[52] (b_vec[52]),     .\b[53] (b_vec[53]),     .\b[54] (b_vec[54]),     .\b[55] (b_vec[55]), 
    .\b[56] (b_vec[56]),     .\b[57] (b_vec[57]),     .\b[58] (b_vec[58]),     .\b[59] (b_vec[59]),     .\b[60] (b_vec[60]),     .\b[61] (b_vec[61]),     .\b[62] (b_vec[62]),     .\b[63] (b_vec[63]), 
    .\b[64] (b_vec[64]),     .\b[65] (b_vec[65]),     .\b[66] (b_vec[66]),     .\b[67] (b_vec[67]),     .\b[68] (b_vec[68]),     .\b[69] (b_vec[69]),     .\b[70] (b_vec[70]),     .\b[71] (b_vec[71]), 
    .\b[72] (b_vec[72]),     .\b[73] (b_vec[73]),     .\b[74] (b_vec[74]),     .\b[75] (b_vec[75]),     .\b[76] (b_vec[76]),     .\b[77] (b_vec[77]),     .\b[78] (b_vec[78]),     .\b[79] (b_vec[79]), 
    .\b[80] (b_vec[80]),     .\b[81] (b_vec[81]),     .\b[82] (b_vec[82]),     .\b[83] (b_vec[83]),     .\b[84] (b_vec[84]),     .\b[85] (b_vec[85]),     .\b[86] (b_vec[86]),     .\b[87] (b_vec[87]), 
    .\b[88] (b_vec[88]),     .\b[89] (b_vec[89]),     .\b[90] (b_vec[90]),     .\b[91] (b_vec[91]),     .\b[92] (b_vec[92]),     .\b[93] (b_vec[93]),     .\b[94] (b_vec[94]),     .\b[95] (b_vec[95]), 
    .\b[96] (b_vec[96]),     .\b[97] (b_vec[97]),     .\b[98] (b_vec[98]),     .\b[99] (b_vec[99]),     .\b[100] (b_vec[100]),     .\b[101] (b_vec[101]),     .\b[102] (b_vec[102]),     .\b[103] (b_vec[103]), 
    .\b[104] (b_vec[104]),     .\b[105] (b_vec[105]),     .\b[106] (b_vec[106]),     .\b[107] (b_vec[107]),     .\b[108] (b_vec[108]),     .\b[109] (b_vec[109]),     .\b[110] (b_vec[110]),     .\b[111] (b_vec[111]), 
    .\b[112] (b_vec[112]),     .\b[113] (b_vec[113]),     .\b[114] (b_vec[114]),     .\b[115] (b_vec[115]),     .\b[116] (b_vec[116]),     .\b[117] (b_vec[117]),     .\b[118] (b_vec[118]),     .\b[119] (b_vec[119]), 
    .\b[120] (b_vec[120]),     .\b[121] (b_vec[121]),     .\b[122] (b_vec[122]),     .\b[123] (b_vec[123]),     .\b[124] (b_vec[124]),     .\b[125] (b_vec[125]),     .\b[126] (b_vec[126]),     .\b[127] (b_vec[127]), 
    .\hypotenuse[0] (hyp_vec[0]),     .\hypotenuse[1] (hyp_vec[1]),     .\hypotenuse[2] (hyp_vec[2]),     .\hypotenuse[3] (hyp_vec[3]),     .\hypotenuse[4] (hyp_vec[4]),     .\hypotenuse[5] (hyp_vec[5]),     .\hypotenuse[6] (hyp_vec[6]),     .\hypotenuse[7] (hyp_vec[7]), 
    .\hypotenuse[8] (hyp_vec[8]),     .\hypotenuse[9] (hyp_vec[9]),     .\hypotenuse[10] (hyp_vec[10]),     .\hypotenuse[11] (hyp_vec[11]),     .\hypotenuse[12] (hyp_vec[12]),     .\hypotenuse[13] (hyp_vec[13]),     .\hypotenuse[14] (hyp_vec[14]),     .\hypotenuse[15] (hyp_vec[15]), 
    .\hypotenuse[16] (hyp_vec[16]),     .\hypotenuse[17] (hyp_vec[17]),     .\hypotenuse[18] (hyp_vec[18]),     .\hypotenuse[19] (hyp_vec[19]),     .\hypotenuse[20] (hyp_vec[20]),     .\hypotenuse[21] (hyp_vec[21]),     .\hypotenuse[22] (hyp_vec[22]),     .\hypotenuse[23] (hyp_vec[23]), 
    .\hypotenuse[24] (hyp_vec[24]),     .\hypotenuse[25] (hyp_vec[25]),     .\hypotenuse[26] (hyp_vec[26]),     .\hypotenuse[27] (hyp_vec[27]),     .\hypotenuse[28] (hyp_vec[28]),     .\hypotenuse[29] (hyp_vec[29]),     .\hypotenuse[30] (hyp_vec[30]),     .\hypotenuse[31] (hyp_vec[31]), 
    .\hypotenuse[32] (hyp_vec[32]),     .\hypotenuse[33] (hyp_vec[33]),     .\hypotenuse[34] (hyp_vec[34]),     .\hypotenuse[35] (hyp_vec[35]),     .\hypotenuse[36] (hyp_vec[36]),     .\hypotenuse[37] (hyp_vec[37]),     .\hypotenuse[38] (hyp_vec[38]),     .\hypotenuse[39] (hyp_vec[39]), 
    .\hypotenuse[40] (hyp_vec[40]),     .\hypotenuse[41] (hyp_vec[41]),     .\hypotenuse[42] (hyp_vec[42]),     .\hypotenuse[43] (hyp_vec[43]),     .\hypotenuse[44] (hyp_vec[44]),     .\hypotenuse[45] (hyp_vec[45]),     .\hypotenuse[46] (hyp_vec[46]),     .\hypotenuse[47] (hyp_vec[47]), 
    .\hypotenuse[48] (hyp_vec[48]),     .\hypotenuse[49] (hyp_vec[49]),     .\hypotenuse[50] (hyp_vec[50]),     .\hypotenuse[51] (hyp_vec[51]),     .\hypotenuse[52] (hyp_vec[52]),     .\hypotenuse[53] (hyp_vec[53]),     .\hypotenuse[54] (hyp_vec[54]),     .\hypotenuse[55] (hyp_vec[55]), 
    .\hypotenuse[56] (hyp_vec[56]),     .\hypotenuse[57] (hyp_vec[57]),     .\hypotenuse[58] (hyp_vec[58]),     .\hypotenuse[59] (hyp_vec[59]),     .\hypotenuse[60] (hyp_vec[60]),     .\hypotenuse[61] (hyp_vec[61]),     .\hypotenuse[62] (hyp_vec[62]),     .\hypotenuse[63] (hyp_vec[63]), 
    .\hypotenuse[64] (hyp_vec[64]),     .\hypotenuse[65] (hyp_vec[65]),     .\hypotenuse[66] (hyp_vec[66]),     .\hypotenuse[67] (hyp_vec[67]),     .\hypotenuse[68] (hyp_vec[68]),     .\hypotenuse[69] (hyp_vec[69]),     .\hypotenuse[70] (hyp_vec[70]),     .\hypotenuse[71] (hyp_vec[71]), 
    .\hypotenuse[72] (hyp_vec[72]),     .\hypotenuse[73] (hyp_vec[73]),     .\hypotenuse[74] (hyp_vec[74]),     .\hypotenuse[75] (hyp_vec[75]),     .\hypotenuse[76] (hyp_vec[76]),     .\hypotenuse[77] (hyp_vec[77]),     .\hypotenuse[78] (hyp_vec[78]),     .\hypotenuse[79] (hyp_vec[79]), 
    .\hypotenuse[80] (hyp_vec[80]),     .\hypotenuse[81] (hyp_vec[81]),     .\hypotenuse[82] (hyp_vec[82]),     .\hypotenuse[83] (hyp_vec[83]),     .\hypotenuse[84] (hyp_vec[84]),     .\hypotenuse[85] (hyp_vec[85]),     .\hypotenuse[86] (hyp_vec[86]),     .\hypotenuse[87] (hyp_vec[87]), 
    .\hypotenuse[88] (hyp_vec[88]),     .\hypotenuse[89] (hyp_vec[89]),     .\hypotenuse[90] (hyp_vec[90]),     .\hypotenuse[91] (hyp_vec[91]),     .\hypotenuse[92] (hyp_vec[92]),     .\hypotenuse[93] (hyp_vec[93]),     .\hypotenuse[94] (hyp_vec[94]),     .\hypotenuse[95] (hyp_vec[95]), 
    .\hypotenuse[96] (hyp_vec[96]),     .\hypotenuse[97] (hyp_vec[97]),     .\hypotenuse[98] (hyp_vec[98]),     .\hypotenuse[99] (hyp_vec[99]),     .\hypotenuse[100] (hyp_vec[100]),     .\hypotenuse[101] (hyp_vec[101]),     .\hypotenuse[102] (hyp_vec[102]),     .\hypotenuse[103] (hyp_vec[103]), 
    .\hypotenuse[104] (hyp_vec[104]),     .\hypotenuse[105] (hyp_vec[105]),     .\hypotenuse[106] (hyp_vec[106]),     .\hypotenuse[107] (hyp_vec[107]),     .\hypotenuse[108] (hyp_vec[108]),     .\hypotenuse[109] (hyp_vec[109]),     .\hypotenuse[110] (hyp_vec[110]),     .\hypotenuse[111] (hyp_vec[111]), 
    .\hypotenuse[112] (hyp_vec[112]),     .\hypotenuse[113] (hyp_vec[113]),     .\hypotenuse[114] (hyp_vec[114]),     .\hypotenuse[115] (hyp_vec[115]),     .\hypotenuse[116] (hyp_vec[116]),     .\hypotenuse[117] (hyp_vec[117]),     .\hypotenuse[118] (hyp_vec[118]),     .\hypotenuse[119] (hyp_vec[119]), 
    .\hypotenuse[120] (hyp_vec[120]),     .\hypotenuse[121] (hyp_vec[121]),     .\hypotenuse[122] (hyp_vec[122]),     .\hypotenuse[123] (hyp_vec[123]),     .\hypotenuse[124] (hyp_vec[124]),     .\hypotenuse[125] (hyp_vec[125]),     .\hypotenuse[126] (hyp_vec[126]),     .\hypotenuse[127] (hyp_vec[127]) 
  );

  integer i;
  parameter STEPS = 64;

  initial begin
    a_vec = 128'b0;
    b_vec = 128'b0;

    #10;

    for (i = 0; i < STEPS; i = i + 1) begin
        if ((i % 2) == 0) a_vec[112] = (i/2 + 0) % 2;
        if ((i % 3) == 0) b_vec[112] = (i/3 + 0 + 1) % 2;
        if ((i % 2) == 0) a_vec[113] = (i/2 + 1) % 2;
        if ((i % 3) == 0) b_vec[113] = (i/3 + 1 + 1) % 2;
        if ((i % 2) == 0) a_vec[114] = (i/2 + 2) % 2;
        if ((i % 3) == 0) b_vec[114] = (i/3 + 2 + 1) % 2;
        if ((i % 2) == 0) a_vec[115] = (i/2 + 3) % 2;
        if ((i % 3) == 0) b_vec[115] = (i/3 + 3 + 1) % 2;
        if ((i % 2) == 0) a_vec[116] = (i/2 + 4) % 2;
        if ((i % 3) == 0) b_vec[116] = (i/3 + 4 + 1) % 2;
        if ((i % 2) == 0) a_vec[117] = (i/2 + 5) % 2;
        if ((i % 3) == 0) b_vec[117] = (i/3 + 5 + 1) % 2;
        if ((i % 2) == 0) a_vec[118] = (i/2 + 6) % 2;
        if ((i % 3) == 0) b_vec[118] = (i/3 + 6 + 1) % 2;
        if ((i % 2) == 0) a_vec[119] = (i/2 + 7) % 2;
        if ((i % 3) == 0) b_vec[119] = (i/3 + 7 + 1) % 2;
        if ((i % 2) == 0) a_vec[120] = (i/2 + 8) % 2;
        if ((i % 3) == 0) b_vec[120] = (i/3 + 8 + 1) % 2;
        if ((i % 2) == 0) a_vec[121] = (i/2 + 9) % 2;
        if ((i % 3) == 0) b_vec[121] = (i/3 + 9 + 1) % 2;
        if ((i % 2) == 0) a_vec[122] = (i/2 + 10) % 2;
        if ((i % 3) == 0) b_vec[122] = (i/3 + 10 + 1) % 2;
        if ((i % 2) == 0) a_vec[123] = (i/2 + 11) % 2;
        if ((i % 3) == 0) b_vec[123] = (i/3 + 11 + 1) % 2;
        if ((i % 2) == 0) a_vec[124] = (i/2 + 12) % 2;
        if ((i % 3) == 0) b_vec[124] = (i/3 + 12 + 1) % 2;
        if ((i % 2) == 0) a_vec[125] = (i/2 + 13) % 2;
        if ((i % 3) == 0) b_vec[125] = (i/3 + 13 + 1) % 2;
        if ((i % 2) == 0) a_vec[126] = (i/2 + 14) % 2;
        if ((i % 3) == 0) b_vec[126] = (i/3 + 14 + 1) % 2;
        if ((i % 2) == 0) a_vec[127] = (i/2 + 15) % 2;
        if ((i % 3) == 0) b_vec[127] = (i/3 + 15 + 1) % 2;
        if ((i % 64) == 0) begin
          a_vec[0] = (i/64 + 0) % 2;
          b_vec[0] = (i/64 + 0 + 1) % 2;
        end
        if ((i % 64) == 0) begin
          a_vec[1] = (i/64 + 1) % 2;
          b_vec[1] = (i/64 + 1 + 1) % 2;
        end
        if ((i % 64) == 0) begin
          a_vec[2] = (i/64 + 2) % 2;
          b_vec[2] = (i/64 + 2 + 1) % 2;
        end
        if ((i % 64) == 0) begin
          a_vec[3] = (i/64 + 3) % 2;
          b_vec[3] = (i/64 + 3 + 1) % 2;
        end
        if ((i % 64) == 0) begin
          a_vec[4] = (i/64 + 4) % 2;
          b_vec[4] = (i/64 + 4 + 1) % 2;
        end
        if ((i % 64) == 0) begin
          a_vec[5] = (i/64 + 5) % 2;
          b_vec[5] = (i/64 + 5 + 1) % 2;
        end
        if ((i % 64) == 0) begin
          a_vec[6] = (i/64 + 6) % 2;
          b_vec[6] = (i/64 + 6 + 1) % 2;
        end
        if ((i % 64) == 0) begin
          a_vec[7] = (i/64 + 7) % 2;
          b_vec[7] = (i/64 + 7 + 1) % 2;
        end

      #1;
      $display("o_sum=%06x", {hyp_vec[0] , hyp_vec[1] , hyp_vec[10] , hyp_vec[100] , hyp_vec[101] , hyp_vec[102] , hyp_vec[103] , hyp_vec[104] , hyp_vec[105] , hyp_vec[106] , hyp_vec[107] , hyp_vec[108] , hyp_vec[109] , hyp_vec[11] , hyp_vec[110] , hyp_vec[111] , hyp_vec[112] , hyp_vec[113] , hyp_vec[114] , hyp_vec[115] , hyp_vec[116] , hyp_vec[117] , hyp_vec[118] , hyp_vec[119] , hyp_vec[12] , hyp_vec[120] , hyp_vec[121] , hyp_vec[122] , hyp_vec[123] , hyp_vec[124] , hyp_vec[125] , hyp_vec[126] , hyp_vec[127] , hyp_vec[13] , hyp_vec[14] , hyp_vec[15] , hyp_vec[16] , hyp_vec[17] , hyp_vec[18] , hyp_vec[19] , hyp_vec[2] , hyp_vec[20] , hyp_vec[21] , hyp_vec[22] , hyp_vec[23] , hyp_vec[24] , hyp_vec[25] , hyp_vec[26] , hyp_vec[27] , hyp_vec[28] , hyp_vec[29] , hyp_vec[3] , hyp_vec[30] , hyp_vec[31] , hyp_vec[32] , hyp_vec[33] , hyp_vec[34] , hyp_vec[35] , hyp_vec[36] , hyp_vec[37] , hyp_vec[38] , hyp_vec[39] , hyp_vec[4] , hyp_vec[40] , hyp_vec[41] , hyp_vec[42] , hyp_vec[43] , hyp_vec[44] , hyp_vec[45] , hyp_vec[46] , hyp_vec[47] , hyp_vec[48] , hyp_vec[49] , hyp_vec[5] , hyp_vec[50] , hyp_vec[51] , hyp_vec[52] , hyp_vec[53] , hyp_vec[54] , hyp_vec[55] , hyp_vec[56] , hyp_vec[57] , hyp_vec[58] , hyp_vec[59] , hyp_vec[6] , hyp_vec[60] , hyp_vec[61] , hyp_vec[62] , hyp_vec[63] , hyp_vec[64] , hyp_vec[65] , hyp_vec[66] , hyp_vec[67] , hyp_vec[68] , hyp_vec[69] , hyp_vec[7] , hyp_vec[70] , hyp_vec[71] , hyp_vec[72] , hyp_vec[73] , hyp_vec[74] , hyp_vec[75] , hyp_vec[76] , hyp_vec[77] , hyp_vec[78] , hyp_vec[79] , hyp_vec[8] , hyp_vec[80] , hyp_vec[81] , hyp_vec[82] , hyp_vec[83] , hyp_vec[84] , hyp_vec[85] , hyp_vec[86] , hyp_vec[87] , hyp_vec[88] , hyp_vec[89] , hyp_vec[9] , hyp_vec[90] , hyp_vec[91] , hyp_vec[92] , hyp_vec[93] , hyp_vec[94] , hyp_vec[95] , hyp_vec[96] , hyp_vec[97] , hyp_vec[98] , hyp_vec[99]});
    end
    $finish;
  end

endmodule
