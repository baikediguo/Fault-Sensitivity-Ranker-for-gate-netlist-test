`timescale 1ns / 1ps

module tb;

  reg pi0000;
  reg pi0001;
  reg pi0002;
  reg pi0003;
  reg pi0004;
  reg pi0005;
  reg pi0006;
  reg pi0007;
  reg pi0008;
  reg pi0009;
  reg pi0010;
  reg pi0011;
  reg pi0012;
  reg pi0013;
  reg pi0014;
  reg pi0015;
  reg pi0016;
  reg pi0017;
  reg pi0018;
  reg pi0019;
  reg pi0020;
  reg pi0021;
  reg pi0022;
  reg pi0023;
  reg pi0024;
  reg pi0025;
  reg pi0026;
  reg pi0027;
  reg pi0028;
  reg pi0029;
  reg pi0030;
  reg pi0031;
  reg pi0032;
  reg pi0033;
  reg pi0034;
  reg pi0035;
  reg pi0036;
  reg pi0037;
  reg pi0038;
  reg pi0039;
  reg pi0040;
  reg pi0041;
  reg pi0042;
  reg pi0043;
  reg pi0044;
  reg pi0045;
  reg pi0046;
  reg pi0047;
  reg pi0048;
  reg pi0049;
  reg pi0050;
  reg pi0051;
  reg pi0052;
  reg pi0053;
  reg pi0054;
  reg pi0055;
  reg pi0056;
  reg pi0057;
  reg pi0058;
  reg pi0059;
  reg pi0060;
  reg pi0061;
  reg pi0062;
  reg pi0063;
  reg pi0064;
  reg pi0065;
  reg pi0066;
  reg pi0067;
  reg pi0068;
  reg pi0069;
  reg pi0070;
  reg pi0071;
  reg pi0072;
  reg pi0073;
  reg pi0074;
  reg pi0075;
  reg pi0076;
  reg pi0077;
  reg pi0078;
  reg pi0079;
  reg pi0080;
  reg pi0081;
  reg pi0082;
  reg pi0083;
  reg pi0084;
  reg pi0085;
  reg pi0086;
  reg pi0087;
  reg pi0088;
  reg pi0089;
  reg pi0090;
  reg pi0091;
  reg pi0092;
  reg pi0093;
  reg pi0094;
  reg pi0095;
  reg pi0096;
  reg pi0097;
  reg pi0098;
  reg pi0099;
  reg pi0100;
  reg pi0101;
  reg pi0102;
  reg pi0103;
  reg pi0104;
  reg pi0105;
  reg pi0106;
  reg pi0107;
  reg pi0108;
  reg pi0109;
  reg pi0110;
  reg pi0111;
  reg pi0112;
  reg pi0113;
  reg pi0114;
  reg pi0115;
  reg pi0116;
  reg pi0117;
  reg pi0118;
  reg pi0119;
  reg pi0120;
  reg pi0121;
  reg pi0122;
  reg pi0123;
  reg pi0124;
  reg pi0125;
  reg pi0126;
  reg pi0127;
  reg pi0128;
  reg pi0129;
  reg pi0130;
  reg pi0131;
  reg pi0132;
  reg pi0133;
  reg pi0134;
  reg pi0135;
  reg pi0136;
  reg pi0137;
  reg pi0138;
  reg pi0139;
  reg pi0140;
  reg pi0141;
  reg pi0142;
  reg pi0143;
  reg pi0144;
  reg pi0145;
  reg pi0146;
  reg pi0147;
  reg pi0148;
  reg pi0149;
  reg pi0150;
  reg pi0151;
  reg pi0152;
  reg pi0153;
  reg pi0154;
  reg pi0155;
  reg pi0156;
  reg pi0157;
  reg pi0158;
  reg pi0159;
  reg pi0160;
  reg pi0161;
  reg pi0162;
  reg pi0163;
  reg pi0164;
  reg pi0165;
  reg pi0166;
  reg pi0167;
  reg pi0168;
  reg pi0169;
  reg pi0170;
  reg pi0171;
  reg pi0172;
  reg pi0173;
  reg pi0174;
  reg pi0175;
  reg pi0176;
  reg pi0177;
  reg pi0178;
  reg pi0179;
  reg pi0180;
  reg pi0181;
  reg pi0182;
  reg pi0183;
  reg pi0184;
  reg pi0185;
  reg pi0186;
  reg pi0187;
  reg pi0188;
  reg pi0189;
  reg pi0190;
  reg pi0191;
  reg pi0192;
  reg pi0193;
  reg pi0194;
  reg pi0195;
  reg pi0196;
  reg pi0197;
  reg pi0198;
  reg pi0199;
  reg pi0200;
  reg pi0201;
  reg pi0202;
  reg pi0203;
  reg pi0204;
  reg pi0205;
  reg pi0206;
  reg pi0207;
  reg pi0208;
  reg pi0209;
  reg pi0210;
  reg pi0211;
  reg pi0212;
  reg pi0213;
  reg pi0214;
  reg pi0215;
  reg pi0216;
  reg pi0217;
  reg pi0218;
  reg pi0219;
  reg pi0220;
  reg pi0221;
  reg pi0222;
  reg pi0223;
  reg pi0224;
  reg pi0225;
  reg pi0226;
  reg pi0227;
  reg pi0228;
  reg pi0229;
  reg pi0230;
  reg pi0231;
  reg pi0232;
  reg pi0233;
  reg pi0234;
  reg pi0235;
  reg pi0236;
  reg pi0237;
  reg pi0238;
  reg pi0239;
  reg pi0240;
  reg pi0241;
  reg pi0242;
  reg pi0243;
  reg pi0244;
  reg pi0245;
  reg pi0246;
  reg pi0247;
  reg pi0248;
  reg pi0249;
  reg pi0250;
  reg pi0251;
  reg pi0252;
  reg pi0253;
  reg pi0254;
  reg pi0255;
  reg pi0256;
  reg pi0257;
  reg pi0258;
  reg pi0259;
  reg pi0260;
  reg pi0261;
  reg pi0262;
  reg pi0263;
  reg pi0264;
  reg pi0265;
  reg pi0266;
  reg pi0267;
  reg pi0268;
  reg pi0269;
  reg pi0270;
  reg pi0271;
  reg pi0272;
  reg pi0273;
  reg pi0274;
  reg pi0275;
  reg pi0276;
  reg pi0277;
  reg pi0278;
  reg pi0279;
  reg pi0280;
  reg pi0281;
  reg pi0282;
  reg pi0283;
  reg pi0284;
  reg pi0285;
  reg pi0286;
  reg pi0287;
  reg pi0288;
  reg pi0289;
  reg pi0290;
  reg pi0291;
  reg pi0292;
  reg pi0293;
  reg pi0294;
  reg pi0295;
  reg pi0296;
  reg pi0297;
  reg pi0298;
  reg pi0299;
  reg pi0300;
  reg pi0301;
  reg pi0302;
  reg pi0303;
  reg pi0304;
  reg pi0305;
  reg pi0306;
  reg pi0307;
  reg pi0308;
  reg pi0309;
  reg pi0310;
  reg pi0311;
  reg pi0312;
  reg pi0313;
  reg pi0314;
  reg pi0315;
  reg pi0316;
  reg pi0317;
  reg pi0318;
  reg pi0319;
  reg pi0320;
  reg pi0321;
  reg pi0322;
  reg pi0323;
  reg pi0324;
  reg pi0325;
  reg pi0326;
  reg pi0327;
  reg pi0328;
  reg pi0329;
  reg pi0330;
  reg pi0331;
  reg pi0332;
  reg pi0333;
  reg pi0334;
  reg pi0335;
  reg pi0336;
  reg pi0337;
  reg pi0338;
  reg pi0339;
  reg pi0340;
  reg pi0341;
  reg pi0342;
  reg pi0343;
  reg pi0344;
  reg pi0345;
  reg pi0346;
  reg pi0347;
  reg pi0348;
  reg pi0349;
  reg pi0350;
  reg pi0351;
  reg pi0352;
  reg pi0353;
  reg pi0354;
  reg pi0355;
  reg pi0356;
  reg pi0357;
  reg pi0358;
  reg pi0359;
  reg pi0360;
  reg pi0361;
  reg pi0362;
  reg pi0363;
  reg pi0364;
  reg pi0365;
  reg pi0366;
  reg pi0367;
  reg pi0368;
  reg pi0369;
  reg pi0370;
  reg pi0371;
  reg pi0372;
  reg pi0373;
  reg pi0374;
  reg pi0375;
  reg pi0376;
  reg pi0377;
  reg pi0378;
  reg pi0379;
  reg pi0380;
  reg pi0381;
  reg pi0382;
  reg pi0383;
  reg pi0384;
  reg pi0385;
  reg pi0386;
  reg pi0387;
  reg pi0388;
  reg pi0389;
  reg pi0390;
  reg pi0391;
  reg pi0392;
  reg pi0393;
  reg pi0394;
  reg pi0395;
  reg pi0396;
  reg pi0397;
  reg pi0398;
  reg pi0399;
  reg pi0400;
  reg pi0401;
  reg pi0402;
  reg pi0403;
  reg pi0404;
  reg pi0405;
  reg pi0406;
  reg pi0407;
  reg pi0408;
  reg pi0409;
  reg pi0410;
  reg pi0411;
  reg pi0412;
  reg pi0413;
  reg pi0414;
  reg pi0415;
  reg pi0416;
  reg pi0417;
  reg pi0418;
  reg pi0419;
  reg pi0420;
  reg pi0421;
  reg pi0422;
  reg pi0423;
  reg pi0424;
  reg pi0425;
  reg pi0426;
  reg pi0427;
  reg pi0428;
  reg pi0429;
  reg pi0430;
  reg pi0431;
  reg pi0432;
  reg pi0433;
  reg pi0434;
  reg pi0435;
  reg pi0436;
  reg pi0437;
  reg pi0438;
  reg pi0439;
  reg pi0440;
  reg pi0441;
  reg pi0442;
  reg pi0443;
  reg pi0444;
  reg pi0445;
  reg pi0446;
  reg pi0447;
  reg pi0448;
  reg pi0449;
  reg pi0450;
  reg pi0451;
  reg pi0452;
  reg pi0453;
  reg pi0454;
  reg pi0455;
  reg pi0456;
  reg pi0457;
  reg pi0458;
  reg pi0459;
  reg pi0460;
  reg pi0461;
  reg pi0462;
  reg pi0463;
  reg pi0464;
  reg pi0465;
  reg pi0466;
  reg pi0467;
  reg pi0468;
  reg pi0469;
  reg pi0470;
  reg pi0471;
  reg pi0472;
  reg pi0473;
  reg pi0474;
  reg pi0475;
  reg pi0476;
  reg pi0477;
  reg pi0478;
  reg pi0479;
  reg pi0480;
  reg pi0481;
  reg pi0482;
  reg pi0483;
  reg pi0484;
  reg pi0485;
  reg pi0486;
  reg pi0487;
  reg pi0488;
  reg pi0489;
  reg pi0490;
  reg pi0491;
  reg pi0492;
  reg pi0493;
  reg pi0494;
  reg pi0495;
  reg pi0496;
  reg pi0497;
  reg pi0498;
  reg pi0499;
  reg pi0500;
  reg pi0501;
  reg pi0502;
  reg pi0503;
  reg pi0504;
  reg pi0505;
  reg pi0506;
  reg pi0507;
  reg pi0508;
  reg pi0509;
  reg pi0510;
  reg pi0511;
  reg pi0512;
  reg pi0513;
  reg pi0514;
  reg pi0515;
  reg pi0516;
  reg pi0517;
  reg pi0518;
  reg pi0519;
  reg pi0520;
  reg pi0521;
  reg pi0522;
  reg pi0523;
  reg pi0524;
  reg pi0525;
  reg pi0526;
  reg pi0527;
  reg pi0528;
  reg pi0529;
  reg pi0530;
  reg pi0531;
  reg pi0532;
  reg pi0533;
  reg pi0534;
  reg pi0535;
  reg pi0536;
  reg pi0537;
  reg pi0538;
  reg pi0539;
  reg pi0540;
  reg pi0541;
  reg pi0542;
  reg pi0543;
  reg pi0544;
  reg pi0545;
  reg pi0546;
  reg pi0547;
  reg pi0548;
  reg pi0549;
  reg pi0550;
  reg pi0551;
  reg pi0552;
  reg pi0553;
  reg pi0554;
  reg pi0555;
  reg pi0556;
  reg pi0557;
  reg pi0558;
  reg pi0559;
  reg pi0560;
  reg pi0561;
  reg pi0562;
  reg pi0563;
  reg pi0564;
  reg pi0565;
  reg pi0566;
  reg pi0567;
  reg pi0568;
  reg pi0569;
  reg pi0570;
  reg pi0571;
  reg pi0572;
  reg pi0573;
  reg pi0574;
  reg pi0575;
  reg pi0576;
  reg pi0577;
  reg pi0578;
  reg pi0579;
  reg pi0580;
  reg pi0581;
  reg pi0582;
  reg pi0583;
  reg pi0584;
  reg pi0585;
  reg pi0586;
  reg pi0587;
  reg pi0588;
  reg pi0589;
  reg pi0590;
  reg pi0591;
  reg pi0592;
  reg pi0593;
  reg pi0594;
  reg pi0595;
  reg pi0596;
  reg pi0597;
  reg pi0598;
  reg pi0599;
  reg pi0600;
  reg pi0601;
  reg pi0602;
  reg pi0603;
  reg pi0604;
  reg pi0605;
  reg pi0606;
  reg pi0607;
  reg pi0608;
  reg pi0609;
  reg pi0610;
  reg pi0611;
  reg pi0612;
  reg pi0613;
  reg pi0614;
  reg pi0615;
  reg pi0616;
  reg pi0617;
  reg pi0618;
  reg pi0619;
  reg pi0620;
  reg pi0621;
  reg pi0622;
  reg pi0623;
  reg pi0624;
  reg pi0625;
  reg pi0626;
  reg pi0627;
  reg pi0628;
  reg pi0629;
  reg pi0630;
  reg pi0631;
  reg pi0632;
  reg pi0633;
  reg pi0634;
  reg pi0635;
  reg pi0636;
  reg pi0637;
  reg pi0638;
  reg pi0639;
  reg pi0640;
  reg pi0641;
  reg pi0642;
  reg pi0643;
  reg pi0644;
  reg pi0645;
  reg pi0646;
  reg pi0647;
  reg pi0648;
  reg pi0649;
  reg pi0650;
  reg pi0651;
  reg pi0652;
  reg pi0653;
  reg pi0654;
  reg pi0655;
  reg pi0656;
  reg pi0657;
  reg pi0658;
  reg pi0659;
  reg pi0660;
  reg pi0661;
  reg pi0662;
  reg pi0663;
  reg pi0664;
  reg pi0665;
  reg pi0666;
  reg pi0667;
  reg pi0668;
  reg pi0669;
  reg pi0670;
  reg pi0671;
  reg pi0672;
  reg pi0673;
  reg pi0674;
  reg pi0675;
  reg pi0676;
  reg pi0677;
  reg pi0678;
  reg pi0679;
  reg pi0680;
  reg pi0681;
  reg pi0682;
  reg pi0683;
  reg pi0684;
  reg pi0685;
  reg pi0686;
  reg pi0687;
  reg pi0688;
  reg pi0689;
  reg pi0690;
  reg pi0691;
  reg pi0692;
  reg pi0693;
  reg pi0694;
  reg pi0695;
  reg pi0696;
  reg pi0697;
  reg pi0698;
  reg pi0699;
  reg pi0700;
  reg pi0701;
  reg pi0702;
  reg pi0703;
  reg pi0704;
  reg pi0705;
  reg pi0706;
  reg pi0707;
  reg pi0708;
  reg pi0709;
  reg pi0710;
  reg pi0711;
  reg pi0712;
  reg pi0713;
  reg pi0714;
  reg pi0715;
  reg pi0716;
  reg pi0717;
  reg pi0718;
  reg pi0719;
  reg pi0720;
  reg pi0721;
  reg pi0722;
  reg pi0723;
  reg pi0724;
  reg pi0725;
  reg pi0726;
  reg pi0727;
  reg pi0728;
  reg pi0729;
  reg pi0730;
  reg pi0731;
  reg pi0732;
  reg pi0733;
  reg pi0734;
  reg pi0735;
  reg pi0736;
  reg pi0737;
  reg pi0738;
  reg pi0739;
  reg pi0740;
  reg pi0741;
  reg pi0742;
  reg pi0743;
  reg pi0744;
  reg pi0745;
  reg pi0746;
  reg pi0747;
  reg pi0748;
  reg pi0749;
  reg pi0750;
  reg pi0751;
  reg pi0752;
  reg pi0753;
  reg pi0754;
  reg pi0755;
  reg pi0756;
  reg pi0757;
  reg pi0758;
  reg pi0759;
  reg pi0760;
  reg pi0761;
  reg pi0762;
  reg pi0763;
  reg pi0764;
  reg pi0765;
  reg pi0766;
  reg pi0767;
  reg pi0768;
  reg pi0769;
  reg pi0770;
  reg pi0771;
  reg pi0772;
  reg pi0773;
  reg pi0774;
  reg pi0775;
  reg pi0776;
  reg pi0777;
  reg pi0778;
  reg pi0779;
  reg pi0780;
  reg pi0781;
  reg pi0782;
  reg pi0783;
  reg pi0784;
  reg pi0785;
  reg pi0786;
  reg pi0787;
  reg pi0788;
  reg pi0789;
  reg pi0790;
  reg pi0791;
  reg pi0792;
  reg pi0793;
  reg pi0794;
  reg pi0795;
  reg pi0796;
  reg pi0797;
  reg pi0798;
  reg pi0799;
  reg pi0800;
  reg pi0801;
  reg pi0802;
  reg pi0803;
  reg pi0804;
  reg pi0805;
  reg pi0806;
  reg pi0807;
  reg pi0808;
  reg pi0809;
  reg pi0810;
  reg pi0811;
  reg pi0812;
  reg pi0813;
  reg pi0814;
  reg pi0815;
  reg pi0816;
  reg pi0817;
  reg pi0818;
  reg pi0819;
  reg pi0820;
  reg pi0821;
  reg pi0822;
  reg pi0823;
  reg pi0824;
  reg pi0825;
  reg pi0826;
  reg pi0827;
  reg pi0828;
  reg pi0829;
  reg pi0830;
  reg pi0831;
  reg pi0832;
  reg pi0833;
  reg pi0834;
  reg pi0835;
  reg pi0836;
  reg pi0837;
  reg pi0838;
  reg pi0839;
  reg pi0840;
  reg pi0841;
  reg pi0842;
  reg pi0843;
  reg pi0844;
  reg pi0845;
  reg pi0846;
  reg pi0847;
  reg pi0848;
  reg pi0849;
  reg pi0850;
  reg pi0851;
  reg pi0852;
  reg pi0853;
  reg pi0854;
  reg pi0855;
  reg pi0856;
  reg pi0857;
  reg pi0858;
  reg pi0859;
  reg pi0860;
  reg pi0861;
  reg pi0862;
  reg pi0863;
  reg pi0864;
  reg pi0865;
  reg pi0866;
  reg pi0867;
  reg pi0868;
  reg pi0869;
  reg pi0870;
  reg pi0871;
  reg pi0872;
  reg pi0873;
  reg pi0874;
  reg pi0875;
  reg pi0876;
  reg pi0877;
  reg pi0878;
  reg pi0879;
  reg pi0880;
  reg pi0881;
  reg pi0882;
  reg pi0883;
  reg pi0884;
  reg pi0885;
  reg pi0886;
  reg pi0887;
  reg pi0888;
  reg pi0889;
  reg pi0890;
  reg pi0891;
  reg pi0892;
  reg pi0893;
  reg pi0894;
  reg pi0895;
  reg pi0896;
  reg pi0897;
  reg pi0898;
  reg pi0899;
  reg pi0900;
  reg pi0901;
  reg pi0902;
  reg pi0903;
  reg pi0904;
  reg pi0905;
  reg pi0906;
  reg pi0907;
  reg pi0908;
  reg pi0909;
  reg pi0910;
  reg pi0911;
  reg pi0912;
  reg pi0913;
  reg pi0914;
  reg pi0915;
  reg pi0916;
  reg pi0917;
  reg pi0918;
  reg pi0919;
  reg pi0920;
  reg pi0921;
  reg pi0922;
  reg pi0923;
  reg pi0924;
  reg pi0925;
  reg pi0926;
  reg pi0927;
  reg pi0928;
  reg pi0929;
  reg pi0930;
  reg pi0931;
  reg pi0932;
  reg pi0933;
  reg pi0934;
  reg pi0935;
  reg pi0936;
  reg pi0937;
  reg pi0938;
  reg pi0939;
  reg pi0940;
  reg pi0941;
  reg pi0942;
  reg pi0943;
  reg pi0944;
  reg pi0945;
  reg pi0946;
  reg pi0947;
  reg pi0948;
  reg pi0949;
  reg pi0950;
  reg pi0951;
  reg pi0952;
  reg pi0953;
  reg pi0954;
  reg pi0955;
  reg pi0956;
  reg pi0957;
  reg pi0958;
  reg pi0959;
  reg pi0960;
  reg pi0961;
  reg pi0962;
  reg pi0963;
  reg pi0964;
  reg pi0965;
  reg pi0966;
  reg pi0967;
  reg pi0968;
  reg pi0969;
  reg pi0970;
  reg pi0971;
  reg pi0972;
  reg pi0973;
  reg pi0974;
  reg pi0975;
  reg pi0976;
  reg pi0977;
  reg pi0978;
  reg pi0979;
  reg pi0980;
  reg pi0981;
  reg pi0982;
  reg pi0983;
  reg pi0984;
  reg pi0985;
  reg pi0986;
  reg pi0987;
  reg pi0988;
  reg pi0989;
  reg pi0990;
  reg pi0991;
  reg pi0992;
  reg pi0993;
  reg pi0994;
  reg pi0995;
  reg pi0996;
  reg pi0997;
  reg pi0998;
  reg pi0999;
  reg pi1000;
  reg pi1001;
  reg pi1002;
  reg pi1003;
  reg pi1004;
  reg pi1005;
  reg pi1006;
  reg pi1007;
  reg pi1008;
  reg pi1009;
  reg pi1010;
  reg pi1011;
  reg pi1012;
  reg pi1013;
  reg pi1014;
  reg pi1015;
  reg pi1016;
  reg pi1017;
  reg pi1018;
  reg pi1019;
  reg pi1020;
  reg pi1021;
  reg pi1022;
  reg pi1023;
  reg pi1024;
  reg pi1025;
  reg pi1026;
  reg pi1027;
  reg pi1028;
  reg pi1029;
  reg pi1030;
  reg pi1031;
  reg pi1032;
  reg pi1033;
  reg pi1034;
  reg pi1035;
  reg pi1036;
  reg pi1037;
  reg pi1038;
  reg pi1039;
  reg pi1040;
  reg pi1041;
  reg pi1042;
  reg pi1043;
  reg pi1044;
  reg pi1045;
  reg pi1046;
  reg pi1047;
  reg pi1048;
  reg pi1049;
  reg pi1050;
  reg pi1051;
  reg pi1052;
  reg pi1053;
  reg pi1054;
  reg pi1055;
  reg pi1056;
  reg pi1057;
  reg pi1058;
  reg pi1059;
  reg pi1060;
  reg pi1061;
  reg pi1062;
  reg pi1063;
  reg pi1064;
  reg pi1065;
  reg pi1066;
  reg pi1067;
  reg pi1068;
  reg pi1069;
  reg pi1070;
  reg pi1071;
  reg pi1072;
  reg pi1073;
  reg pi1074;
  reg pi1075;
  reg pi1076;
  reg pi1077;
  reg pi1078;
  reg pi1079;
  reg pi1080;
  reg pi1081;
  reg pi1082;
  reg pi1083;
  reg pi1084;
  reg pi1085;
  reg pi1086;
  reg pi1087;
  reg pi1088;
  reg pi1089;
  reg pi1090;
  reg pi1091;
  reg pi1092;
  reg pi1093;
  reg pi1094;
  reg pi1095;
  reg pi1096;
  reg pi1097;
  reg pi1098;
  reg pi1099;
  reg pi1100;
  reg pi1101;
  reg pi1102;
  reg pi1103;
  reg pi1104;
  reg pi1105;
  reg pi1106;
  reg pi1107;
  reg pi1108;
  reg pi1109;
  reg pi1110;
  reg pi1111;
  reg pi1112;
  reg pi1113;
  reg pi1114;
  reg pi1115;
  reg pi1116;
  reg pi1117;
  reg pi1118;
  reg pi1119;
  reg pi1120;
  reg pi1121;
  reg pi1122;
  reg pi1123;
  reg pi1124;
  reg pi1125;
  reg pi1126;
  reg pi1127;
  reg pi1128;
  reg pi1129;
  reg pi1130;
  reg pi1131;
  reg pi1132;
  reg pi1133;
  reg pi1134;
  reg pi1135;
  reg pi1136;
  reg pi1137;
  reg pi1138;
  reg pi1139;
  reg pi1140;
  reg pi1141;
  reg pi1142;
  reg pi1143;
  reg pi1144;
  reg pi1145;
  reg pi1146;
  reg pi1147;
  reg pi1148;
  reg pi1149;
  reg pi1150;
  reg pi1151;
  reg pi1152;
  reg pi1153;
  reg pi1154;
  reg pi1155;
  reg pi1156;
  reg pi1157;
  reg pi1158;
  reg pi1159;
  reg pi1160;
  reg pi1161;
  reg pi1162;
  reg pi1163;
  reg pi1164;
  reg pi1165;
  reg pi1166;
  reg pi1167;
  reg pi1168;
  reg pi1169;
  reg pi1170;
  reg pi1171;
  reg pi1172;
  reg pi1173;
  reg pi1174;
  reg pi1175;
  reg pi1176;
  reg pi1177;
  reg pi1178;
  reg pi1179;
  reg pi1180;
  reg pi1181;
  reg pi1182;
  reg pi1183;
  reg pi1184;
  reg pi1185;
  reg pi1186;
  reg pi1187;
  reg pi1188;
  reg pi1189;
  reg pi1190;
  reg pi1191;
  reg pi1192;
  reg pi1193;
  reg pi1194;
  reg pi1195;
  reg pi1196;
  reg pi1197;
  reg pi1198;
  reg pi1199;
  reg pi1200;
  reg pi1201;
  reg pi1202;
  reg pi1203;
  wire po0000;
  wire po0001;
  wire po0002;
  wire po0003;
  wire po0004;
  wire po0005;
  wire po0006;
  wire po0007;
  wire po0008;
  wire po0009;
  wire po0010;
  wire po0011;
  wire po0012;
  wire po0013;
  wire po0014;
  wire po0015;
  wire po0016;
  wire po0017;
  wire po0018;
  wire po0019;
  wire po0020;
  wire po0021;
  wire po0022;
  wire po0023;
  wire po0024;
  wire po0025;
  wire po0026;
  wire po0027;
  wire po0028;
  wire po0029;
  wire po0030;
  wire po0031;
  wire po0032;
  wire po0033;
  wire po0034;
  wire po0035;
  wire po0036;
  wire po0037;
  wire po0038;
  wire po0039;
  wire po0040;
  wire po0041;
  wire po0042;
  wire po0043;
  wire po0044;
  wire po0045;
  wire po0046;
  wire po0047;
  wire po0048;
  wire po0049;
  wire po0050;
  wire po0051;
  wire po0052;
  wire po0053;
  wire po0054;
  wire po0055;
  wire po0056;
  wire po0057;
  wire po0058;
  wire po0059;
  wire po0060;
  wire po0061;
  wire po0062;
  wire po0063;
  wire po0064;
  wire po0065;
  wire po0066;
  wire po0067;
  wire po0068;
  wire po0069;
  wire po0070;
  wire po0071;
  wire po0072;
  wire po0073;
  wire po0074;
  wire po0075;
  wire po0076;
  wire po0077;
  wire po0078;
  wire po0079;
  wire po0080;
  wire po0081;
  wire po0082;
  wire po0083;
  wire po0084;
  wire po0085;
  wire po0086;
  wire po0087;
  wire po0088;
  wire po0089;
  wire po0090;
  wire po0091;
  wire po0092;
  wire po0093;
  wire po0094;
  wire po0095;
  wire po0096;
  wire po0097;
  wire po0098;
  wire po0099;
  wire po0100;
  wire po0101;
  wire po0102;
  wire po0103;
  wire po0104;
  wire po0105;
  wire po0106;
  wire po0107;
  wire po0108;
  wire po0109;
  wire po0110;
  wire po0111;
  wire po0112;
  wire po0113;
  wire po0114;
  wire po0115;
  wire po0116;
  wire po0117;
  wire po0118;
  wire po0119;
  wire po0120;
  wire po0121;
  wire po0122;
  wire po0123;
  wire po0124;
  wire po0125;
  wire po0126;
  wire po0127;
  wire po0128;
  wire po0129;
  wire po0130;
  wire po0131;
  wire po0132;
  wire po0133;
  wire po0134;
  wire po0135;
  wire po0136;
  wire po0137;
  wire po0138;
  wire po0139;
  wire po0140;
  wire po0141;
  wire po0142;
  wire po0143;
  wire po0144;
  wire po0145;
  wire po0146;
  wire po0147;
  wire po0148;
  wire po0149;
  wire po0150;
  wire po0151;
  wire po0152;
  wire po0153;
  wire po0154;
  wire po0155;
  wire po0156;
  wire po0157;
  wire po0158;
  wire po0159;
  wire po0160;
  wire po0161;
  wire po0162;
  wire po0163;
  wire po0164;
  wire po0165;
  wire po0166;
  wire po0167;
  wire po0168;
  wire po0169;
  wire po0170;
  wire po0171;
  wire po0172;
  wire po0173;
  wire po0174;
  wire po0175;
  wire po0176;
  wire po0177;
  wire po0178;
  wire po0179;
  wire po0180;
  wire po0181;
  wire po0182;
  wire po0183;
  wire po0184;
  wire po0185;
  wire po0186;
  wire po0187;
  wire po0188;
  wire po0189;
  wire po0190;
  wire po0191;
  wire po0192;
  wire po0193;
  wire po0194;
  wire po0195;
  wire po0196;
  wire po0197;
  wire po0198;
  wire po0199;
  wire po0200;
  wire po0201;
  wire po0202;
  wire po0203;
  wire po0204;
  wire po0205;
  wire po0206;
  wire po0207;
  wire po0208;
  wire po0209;
  wire po0210;
  wire po0211;
  wire po0212;
  wire po0213;
  wire po0214;
  wire po0215;
  wire po0216;
  wire po0217;
  wire po0218;
  wire po0219;
  wire po0220;
  wire po0221;
  wire po0222;
  wire po0223;
  wire po0224;
  wire po0225;
  wire po0226;
  wire po0227;
  wire po0228;
  wire po0229;
  wire po0230;
  wire po0231;
  wire po0232;
  wire po0233;
  wire po0234;
  wire po0235;
  wire po0236;
  wire po0237;
  wire po0238;
  wire po0239;
  wire po0240;
  wire po0241;
  wire po0242;
  wire po0243;
  wire po0244;
  wire po0245;
  wire po0246;
  wire po0247;
  wire po0248;
  wire po0249;
  wire po0250;
  wire po0251;
  wire po0252;
  wire po0253;
  wire po0254;
  wire po0255;
  wire po0256;
  wire po0257;
  wire po0258;
  wire po0259;
  wire po0260;
  wire po0261;
  wire po0262;
  wire po0263;
  wire po0264;
  wire po0265;
  wire po0266;
  wire po0267;
  wire po0268;
  wire po0269;
  wire po0270;
  wire po0271;
  wire po0272;
  wire po0273;
  wire po0274;
  wire po0275;
  wire po0276;
  wire po0277;
  wire po0278;
  wire po0279;
  wire po0280;
  wire po0281;
  wire po0282;
  wire po0283;
  wire po0284;
  wire po0285;
  wire po0286;
  wire po0287;
  wire po0288;
  wire po0289;
  wire po0290;
  wire po0291;
  wire po0292;
  wire po0293;
  wire po0294;
  wire po0295;
  wire po0296;
  wire po0297;
  wire po0298;
  wire po0299;
  wire po0300;
  wire po0301;
  wire po0302;
  wire po0303;
  wire po0304;
  wire po0305;
  wire po0306;
  wire po0307;
  wire po0308;
  wire po0309;
  wire po0310;
  wire po0311;
  wire po0312;
  wire po0313;
  wire po0314;
  wire po0315;
  wire po0316;
  wire po0317;
  wire po0318;
  wire po0319;
  wire po0320;
  wire po0321;
  wire po0322;
  wire po0323;
  wire po0324;
  wire po0325;
  wire po0326;
  wire po0327;
  wire po0328;
  wire po0329;
  wire po0330;
  wire po0331;
  wire po0332;
  wire po0333;
  wire po0334;
  wire po0335;
  wire po0336;
  wire po0337;
  wire po0338;
  wire po0339;
  wire po0340;
  wire po0341;
  wire po0342;
  wire po0343;
  wire po0344;
  wire po0345;
  wire po0346;
  wire po0347;
  wire po0348;
  wire po0349;
  wire po0350;
  wire po0351;
  wire po0352;
  wire po0353;
  wire po0354;
  wire po0355;
  wire po0356;
  wire po0357;
  wire po0358;
  wire po0359;
  wire po0360;
  wire po0361;
  wire po0362;
  wire po0363;
  wire po0364;
  wire po0365;
  wire po0366;
  wire po0367;
  wire po0368;
  wire po0369;
  wire po0370;
  wire po0371;
  wire po0372;
  wire po0373;
  wire po0374;
  wire po0375;
  wire po0376;
  wire po0377;
  wire po0378;
  wire po0379;
  wire po0380;
  wire po0381;
  wire po0382;
  wire po0383;
  wire po0384;
  wire po0385;
  wire po0386;
  wire po0387;
  wire po0388;
  wire po0389;
  wire po0390;
  wire po0391;
  wire po0392;
  wire po0393;
  wire po0394;
  wire po0395;
  wire po0396;
  wire po0397;
  wire po0398;
  wire po0399;
  wire po0400;
  wire po0401;
  wire po0402;
  wire po0403;
  wire po0404;
  wire po0405;
  wire po0406;
  wire po0407;
  wire po0408;
  wire po0409;
  wire po0410;
  wire po0411;
  wire po0412;
  wire po0413;
  wire po0414;
  wire po0415;
  wire po0416;
  wire po0417;
  wire po0418;
  wire po0419;
  wire po0420;
  wire po0421;
  wire po0422;
  wire po0423;
  wire po0424;
  wire po0425;
  wire po0426;
  wire po0427;
  wire po0428;
  wire po0429;
  wire po0430;
  wire po0431;
  wire po0432;
  wire po0433;
  wire po0434;
  wire po0435;
  wire po0436;
  wire po0437;
  wire po0438;
  wire po0439;
  wire po0440;
  wire po0441;
  wire po0442;
  wire po0443;
  wire po0444;
  wire po0445;
  wire po0446;
  wire po0447;
  wire po0448;
  wire po0449;
  wire po0450;
  wire po0451;
  wire po0452;
  wire po0453;
  wire po0454;
  wire po0455;
  wire po0456;
  wire po0457;
  wire po0458;
  wire po0459;
  wire po0460;
  wire po0461;
  wire po0462;
  wire po0463;
  wire po0464;
  wire po0465;
  wire po0466;
  wire po0467;
  wire po0468;
  wire po0469;
  wire po0470;
  wire po0471;
  wire po0472;
  wire po0473;
  wire po0474;
  wire po0475;
  wire po0476;
  wire po0477;
  wire po0478;
  wire po0479;
  wire po0480;
  wire po0481;
  wire po0482;
  wire po0483;
  wire po0484;
  wire po0485;
  wire po0486;
  wire po0487;
  wire po0488;
  wire po0489;
  wire po0490;
  wire po0491;
  wire po0492;
  wire po0493;
  wire po0494;
  wire po0495;
  wire po0496;
  wire po0497;
  wire po0498;
  wire po0499;
  wire po0500;
  wire po0501;
  wire po0502;
  wire po0503;
  wire po0504;
  wire po0505;
  wire po0506;
  wire po0507;
  wire po0508;
  wire po0509;
  wire po0510;
  wire po0511;
  wire po0512;
  wire po0513;
  wire po0514;
  wire po0515;
  wire po0516;
  wire po0517;
  wire po0518;
  wire po0519;
  wire po0520;
  wire po0521;
  wire po0522;
  wire po0523;
  wire po0524;
  wire po0525;
  wire po0526;
  wire po0527;
  wire po0528;
  wire po0529;
  wire po0530;
  wire po0531;
  wire po0532;
  wire po0533;
  wire po0534;
  wire po0535;
  wire po0536;
  wire po0537;
  wire po0538;
  wire po0539;
  wire po0540;
  wire po0541;
  wire po0542;
  wire po0543;
  wire po0544;
  wire po0545;
  wire po0546;
  wire po0547;
  wire po0548;
  wire po0549;
  wire po0550;
  wire po0551;
  wire po0552;
  wire po0553;
  wire po0554;
  wire po0555;
  wire po0556;
  wire po0557;
  wire po0558;
  wire po0559;
  wire po0560;
  wire po0561;
  wire po0562;
  wire po0563;
  wire po0564;
  wire po0565;
  wire po0566;
  wire po0567;
  wire po0568;
  wire po0569;
  wire po0570;
  wire po0571;
  wire po0572;
  wire po0573;
  wire po0574;
  wire po0575;
  wire po0576;
  wire po0577;
  wire po0578;
  wire po0579;
  wire po0580;
  wire po0581;
  wire po0582;
  wire po0583;
  wire po0584;
  wire po0585;
  wire po0586;
  wire po0587;
  wire po0588;
  wire po0589;
  wire po0590;
  wire po0591;
  wire po0592;
  wire po0593;
  wire po0594;
  wire po0595;
  wire po0596;
  wire po0597;
  wire po0598;
  wire po0599;
  wire po0600;
  wire po0601;
  wire po0602;
  wire po0603;
  wire po0604;
  wire po0605;
  wire po0606;
  wire po0607;
  wire po0608;
  wire po0609;
  wire po0610;
  wire po0611;
  wire po0612;
  wire po0613;
  wire po0614;
  wire po0615;
  wire po0616;
  wire po0617;
  wire po0618;
  wire po0619;
  wire po0620;
  wire po0621;
  wire po0622;
  wire po0623;
  wire po0624;
  wire po0625;
  wire po0626;
  wire po0627;
  wire po0628;
  wire po0629;
  wire po0630;
  wire po0631;
  wire po0632;
  wire po0633;
  wire po0634;
  wire po0635;
  wire po0636;
  wire po0637;
  wire po0638;
  wire po0639;
  wire po0640;
  wire po0641;
  wire po0642;
  wire po0643;
  wire po0644;
  wire po0645;
  wire po0646;
  wire po0647;
  wire po0648;
  wire po0649;
  wire po0650;
  wire po0651;
  wire po0652;
  wire po0653;
  wire po0654;
  wire po0655;
  wire po0656;
  wire po0657;
  wire po0658;
  wire po0659;
  wire po0660;
  wire po0661;
  wire po0662;
  wire po0663;
  wire po0664;
  wire po0665;
  wire po0666;
  wire po0667;
  wire po0668;
  wire po0669;
  wire po0670;
  wire po0671;
  wire po0672;
  wire po0673;
  wire po0674;
  wire po0675;
  wire po0676;
  wire po0677;
  wire po0678;
  wire po0679;
  wire po0680;
  wire po0681;
  wire po0682;
  wire po0683;
  wire po0684;
  wire po0685;
  wire po0686;
  wire po0687;
  wire po0688;
  wire po0689;
  wire po0690;
  wire po0691;
  wire po0692;
  wire po0693;
  wire po0694;
  wire po0695;
  wire po0696;
  wire po0697;
  wire po0698;
  wire po0699;
  wire po0700;
  wire po0701;
  wire po0702;
  wire po0703;
  wire po0704;
  wire po0705;
  wire po0706;
  wire po0707;
  wire po0708;
  wire po0709;
  wire po0710;
  wire po0711;
  wire po0712;
  wire po0713;
  wire po0714;
  wire po0715;
  wire po0716;
  wire po0717;
  wire po0718;
  wire po0719;
  wire po0720;
  wire po0721;
  wire po0722;
  wire po0723;
  wire po0724;
  wire po0725;
  wire po0726;
  wire po0727;
  wire po0728;
  wire po0729;
  wire po0730;
  wire po0731;
  wire po0732;
  wire po0733;
  wire po0734;
  wire po0735;
  wire po0736;
  wire po0737;
  wire po0738;
  wire po0739;
  wire po0740;
  wire po0741;
  wire po0742;
  wire po0743;
  wire po0744;
  wire po0745;
  wire po0746;
  wire po0747;
  wire po0748;
  wire po0749;
  wire po0750;
  wire po0751;
  wire po0752;
  wire po0753;
  wire po0754;
  wire po0755;
  wire po0756;
  wire po0757;
  wire po0758;
  wire po0759;
  wire po0760;
  wire po0761;
  wire po0762;
  wire po0763;
  wire po0764;
  wire po0765;
  wire po0766;
  wire po0767;
  wire po0768;
  wire po0769;
  wire po0770;
  wire po0771;
  wire po0772;
  wire po0773;
  wire po0774;
  wire po0775;
  wire po0776;
  wire po0777;
  wire po0778;
  wire po0779;
  wire po0780;
  wire po0781;
  wire po0782;
  wire po0783;
  wire po0784;
  wire po0785;
  wire po0786;
  wire po0787;
  wire po0788;
  wire po0789;
  wire po0790;
  wire po0791;
  wire po0792;
  wire po0793;
  wire po0794;
  wire po0795;
  wire po0796;
  wire po0797;
  wire po0798;
  wire po0799;
  wire po0800;
  wire po0801;
  wire po0802;
  wire po0803;
  wire po0804;
  wire po0805;
  wire po0806;
  wire po0807;
  wire po0808;
  wire po0809;
  wire po0810;
  wire po0811;
  wire po0812;
  wire po0813;
  wire po0814;
  wire po0815;
  wire po0816;
  wire po0817;
  wire po0818;
  wire po0819;
  wire po0820;
  wire po0821;
  wire po0822;
  wire po0823;
  wire po0824;
  wire po0825;
  wire po0826;
  wire po0827;
  wire po0828;
  wire po0829;
  wire po0830;
  wire po0831;
  wire po0832;
  wire po0833;
  wire po0834;
  wire po0835;
  wire po0836;
  wire po0837;
  wire po0838;
  wire po0839;
  wire po0840;
  wire po0841;
  wire po0842;
  wire po0843;
  wire po0844;
  wire po0845;
  wire po0846;
  wire po0847;
  wire po0848;
  wire po0849;
  wire po0850;
  wire po0851;
  wire po0852;
  wire po0853;
  wire po0854;
  wire po0855;
  wire po0856;
  wire po0857;
  wire po0858;
  wire po0859;
  wire po0860;
  wire po0861;
  wire po0862;
  wire po0863;
  wire po0864;
  wire po0865;
  wire po0866;
  wire po0867;
  wire po0868;
  wire po0869;
  wire po0870;
  wire po0871;
  wire po0872;
  wire po0873;
  wire po0874;
  wire po0875;
  wire po0876;
  wire po0877;
  wire po0878;
  wire po0879;
  wire po0880;
  wire po0881;
  wire po0882;
  wire po0883;
  wire po0884;
  wire po0885;
  wire po0886;
  wire po0887;
  wire po0888;
  wire po0889;
  wire po0890;
  wire po0891;
  wire po0892;
  wire po0893;
  wire po0894;
  wire po0895;
  wire po0896;
  wire po0897;
  wire po0898;
  wire po0899;
  wire po0900;
  wire po0901;
  wire po0902;
  wire po0903;
  wire po0904;
  wire po0905;
  wire po0906;
  wire po0907;
  wire po0908;
  wire po0909;
  wire po0910;
  wire po0911;
  wire po0912;
  wire po0913;
  wire po0914;
  wire po0915;
  wire po0916;
  wire po0917;
  wire po0918;
  wire po0919;
  wire po0920;
  wire po0921;
  wire po0922;
  wire po0923;
  wire po0924;
  wire po0925;
  wire po0926;
  wire po0927;
  wire po0928;
  wire po0929;
  wire po0930;
  wire po0931;
  wire po0932;
  wire po0933;
  wire po0934;
  wire po0935;
  wire po0936;
  wire po0937;
  wire po0938;
  wire po0939;
  wire po0940;
  wire po0941;
  wire po0942;
  wire po0943;
  wire po0944;
  wire po0945;
  wire po0946;
  wire po0947;
  wire po0948;
  wire po0949;
  wire po0950;
  wire po0951;
  wire po0952;
  wire po0953;
  wire po0954;
  wire po0955;
  wire po0956;
  wire po0957;
  wire po0958;
  wire po0959;
  wire po0960;
  wire po0961;
  wire po0962;
  wire po0963;
  wire po0964;
  wire po0965;
  wire po0966;
  wire po0967;
  wire po0968;
  wire po0969;
  wire po0970;
  wire po0971;
  wire po0972;
  wire po0973;
  wire po0974;
  wire po0975;
  wire po0976;
  wire po0977;
  wire po0978;
  wire po0979;
  wire po0980;
  wire po0981;
  wire po0982;
  wire po0983;
  wire po0984;
  wire po0985;
  wire po0986;
  wire po0987;
  wire po0988;
  wire po0989;
  wire po0990;
  wire po0991;
  wire po0992;
  wire po0993;
  wire po0994;
  wire po0995;
  wire po0996;
  wire po0997;
  wire po0998;
  wire po0999;
  wire po1000;
  wire po1001;
  wire po1002;
  wire po1003;
  wire po1004;
  wire po1005;
  wire po1006;
  wire po1007;
  wire po1008;
  wire po1009;
  wire po1010;
  wire po1011;
  wire po1012;
  wire po1013;
  wire po1014;
  wire po1015;
  wire po1016;
  wire po1017;
  wire po1018;
  wire po1019;
  wire po1020;
  wire po1021;
  wire po1022;
  wire po1023;
  wire po1024;
  wire po1025;
  wire po1026;
  wire po1027;
  wire po1028;
  wire po1029;
  wire po1030;
  wire po1031;
  wire po1032;
  wire po1033;
  wire po1034;
  wire po1035;
  wire po1036;
  wire po1037;
  wire po1038;
  wire po1039;
  wire po1040;
  wire po1041;
  wire po1042;
  wire po1043;
  wire po1044;
  wire po1045;
  wire po1046;
  wire po1047;
  wire po1048;
  wire po1049;
  wire po1050;
  wire po1051;
  wire po1052;
  wire po1053;
  wire po1054;
  wire po1055;
  wire po1056;
  wire po1057;
  wire po1058;
  wire po1059;
  wire po1060;
  wire po1061;
  wire po1062;
  wire po1063;
  wire po1064;
  wire po1065;
  wire po1066;
  wire po1067;
  wire po1068;
  wire po1069;
  wire po1070;
  wire po1071;
  wire po1072;
  wire po1073;
  wire po1074;
  wire po1075;
  wire po1076;
  wire po1077;
  wire po1078;
  wire po1079;
  wire po1080;
  wire po1081;
  wire po1082;
  wire po1083;
  wire po1084;
  wire po1085;
  wire po1086;
  wire po1087;
  wire po1088;
  wire po1089;
  wire po1090;
  wire po1091;
  wire po1092;
  wire po1093;
  wire po1094;
  wire po1095;
  wire po1096;
  wire po1097;
  wire po1098;
  wire po1099;
  wire po1100;
  wire po1101;
  wire po1102;
  wire po1103;
  wire po1104;
  wire po1105;
  wire po1106;
  wire po1107;
  wire po1108;
  wire po1109;
  wire po1110;
  wire po1111;
  wire po1112;
  wire po1113;
  wire po1114;
  wire po1115;
  wire po1116;
  wire po1117;
  wire po1118;
  wire po1119;
  wire po1120;
  wire po1121;
  wire po1122;
  wire po1123;
  wire po1124;
  wire po1125;
  wire po1126;
  wire po1127;
  wire po1128;
  wire po1129;
  wire po1130;
  wire po1131;
  wire po1132;
  wire po1133;
  wire po1134;
  wire po1135;
  wire po1136;
  wire po1137;
  wire po1138;
  wire po1139;
  wire po1140;
  wire po1141;
  wire po1142;
  wire po1143;
  wire po1144;
  wire po1145;
  wire po1146;
  wire po1147;
  wire po1148;
  wire po1149;
  wire po1150;
  wire po1151;
  wire po1152;
  wire po1153;
  wire po1154;
  wire po1155;
  wire po1156;
  wire po1157;
  wire po1158;
  wire po1159;
  wire po1160;
  wire po1161;
  wire po1162;
  wire po1163;
  wire po1164;
  wire po1165;
  wire po1166;
  wire po1167;
  wire po1168;
  wire po1169;
  wire po1170;
  wire po1171;
  wire po1172;
  wire po1173;
  wire po1174;
  wire po1175;
  wire po1176;
  wire po1177;
  wire po1178;
  wire po1179;
  wire po1180;
  wire po1181;
  wire po1182;
  wire po1183;
  wire po1184;
  wire po1185;
  wire po1186;
  wire po1187;
  wire po1188;
  wire po1189;
  wire po1190;
  wire po1191;
  wire po1192;
  wire po1193;
  wire po1194;
  wire po1195;
  wire po1196;
  wire po1197;
  wire po1198;
  wire po1199;
  wire po1200;
  wire po1201;
  wire po1202;
  wire po1203;
  wire po1204;
  wire po1205;
  wire po1206;
  wire po1207;
  wire po1208;
  wire po1209;
  wire po1210;
  wire po1211;
  wire po1212;
  wire po1213;
  wire po1214;
  wire po1215;
  wire po1216;
  wire po1217;
  wire po1218;
  wire po1219;
  wire po1220;
  wire po1221;
  wire po1222;
  wire po1223;
  wire po1224;
  wire po1225;
  wire po1226;
  wire po1227;
  wire po1228;
  wire po1229;
  wire po1230;

  // DUT (combinational)
  mem_ctrl uut (
    .pi0000(pi0000),
    .pi0001(pi0001),
    .pi0002(pi0002),
    .pi0003(pi0003),
    .pi0004(pi0004),
    .pi0005(pi0005),
    .pi0006(pi0006),
    .pi0007(pi0007),
    .pi0008(pi0008),
    .pi0009(pi0009),
    .pi0010(pi0010),
    .pi0011(pi0011),
    .pi0012(pi0012),
    .pi0013(pi0013),
    .pi0014(pi0014),
    .pi0015(pi0015),
    .pi0016(pi0016),
    .pi0017(pi0017),
    .pi0018(pi0018),
    .pi0019(pi0019),
    .pi0020(pi0020),
    .pi0021(pi0021),
    .pi0022(pi0022),
    .pi0023(pi0023),
    .pi0024(pi0024),
    .pi0025(pi0025),
    .pi0026(pi0026),
    .pi0027(pi0027),
    .pi0028(pi0028),
    .pi0029(pi0029),
    .pi0030(pi0030),
    .pi0031(pi0031),
    .pi0032(pi0032),
    .pi0033(pi0033),
    .pi0034(pi0034),
    .pi0035(pi0035),
    .pi0036(pi0036),
    .pi0037(pi0037),
    .pi0038(pi0038),
    .pi0039(pi0039),
    .pi0040(pi0040),
    .pi0041(pi0041),
    .pi0042(pi0042),
    .pi0043(pi0043),
    .pi0044(pi0044),
    .pi0045(pi0045),
    .pi0046(pi0046),
    .pi0047(pi0047),
    .pi0048(pi0048),
    .pi0049(pi0049),
    .pi0050(pi0050),
    .pi0051(pi0051),
    .pi0052(pi0052),
    .pi0053(pi0053),
    .pi0054(pi0054),
    .pi0055(pi0055),
    .pi0056(pi0056),
    .pi0057(pi0057),
    .pi0058(pi0058),
    .pi0059(pi0059),
    .pi0060(pi0060),
    .pi0061(pi0061),
    .pi0062(pi0062),
    .pi0063(pi0063),
    .pi0064(pi0064),
    .pi0065(pi0065),
    .pi0066(pi0066),
    .pi0067(pi0067),
    .pi0068(pi0068),
    .pi0069(pi0069),
    .pi0070(pi0070),
    .pi0071(pi0071),
    .pi0072(pi0072),
    .pi0073(pi0073),
    .pi0074(pi0074),
    .pi0075(pi0075),
    .pi0076(pi0076),
    .pi0077(pi0077),
    .pi0078(pi0078),
    .pi0079(pi0079),
    .pi0080(pi0080),
    .pi0081(pi0081),
    .pi0082(pi0082),
    .pi0083(pi0083),
    .pi0084(pi0084),
    .pi0085(pi0085),
    .pi0086(pi0086),
    .pi0087(pi0087),
    .pi0088(pi0088),
    .pi0089(pi0089),
    .pi0090(pi0090),
    .pi0091(pi0091),
    .pi0092(pi0092),
    .pi0093(pi0093),
    .pi0094(pi0094),
    .pi0095(pi0095),
    .pi0096(pi0096),
    .pi0097(pi0097),
    .pi0098(pi0098),
    .pi0099(pi0099),
    .pi0100(pi0100),
    .pi0101(pi0101),
    .pi0102(pi0102),
    .pi0103(pi0103),
    .pi0104(pi0104),
    .pi0105(pi0105),
    .pi0106(pi0106),
    .pi0107(pi0107),
    .pi0108(pi0108),
    .pi0109(pi0109),
    .pi0110(pi0110),
    .pi0111(pi0111),
    .pi0112(pi0112),
    .pi0113(pi0113),
    .pi0114(pi0114),
    .pi0115(pi0115),
    .pi0116(pi0116),
    .pi0117(pi0117),
    .pi0118(pi0118),
    .pi0119(pi0119),
    .pi0120(pi0120),
    .pi0121(pi0121),
    .pi0122(pi0122),
    .pi0123(pi0123),
    .pi0124(pi0124),
    .pi0125(pi0125),
    .pi0126(pi0126),
    .pi0127(pi0127),
    .pi0128(pi0128),
    .pi0129(pi0129),
    .pi0130(pi0130),
    .pi0131(pi0131),
    .pi0132(pi0132),
    .pi0133(pi0133),
    .pi0134(pi0134),
    .pi0135(pi0135),
    .pi0136(pi0136),
    .pi0137(pi0137),
    .pi0138(pi0138),
    .pi0139(pi0139),
    .pi0140(pi0140),
    .pi0141(pi0141),
    .pi0142(pi0142),
    .pi0143(pi0143),
    .pi0144(pi0144),
    .pi0145(pi0145),
    .pi0146(pi0146),
    .pi0147(pi0147),
    .pi0148(pi0148),
    .pi0149(pi0149),
    .pi0150(pi0150),
    .pi0151(pi0151),
    .pi0152(pi0152),
    .pi0153(pi0153),
    .pi0154(pi0154),
    .pi0155(pi0155),
    .pi0156(pi0156),
    .pi0157(pi0157),
    .pi0158(pi0158),
    .pi0159(pi0159),
    .pi0160(pi0160),
    .pi0161(pi0161),
    .pi0162(pi0162),
    .pi0163(pi0163),
    .pi0164(pi0164),
    .pi0165(pi0165),
    .pi0166(pi0166),
    .pi0167(pi0167),
    .pi0168(pi0168),
    .pi0169(pi0169),
    .pi0170(pi0170),
    .pi0171(pi0171),
    .pi0172(pi0172),
    .pi0173(pi0173),
    .pi0174(pi0174),
    .pi0175(pi0175),
    .pi0176(pi0176),
    .pi0177(pi0177),
    .pi0178(pi0178),
    .pi0179(pi0179),
    .pi0180(pi0180),
    .pi0181(pi0181),
    .pi0182(pi0182),
    .pi0183(pi0183),
    .pi0184(pi0184),
    .pi0185(pi0185),
    .pi0186(pi0186),
    .pi0187(pi0187),
    .pi0188(pi0188),
    .pi0189(pi0189),
    .pi0190(pi0190),
    .pi0191(pi0191),
    .pi0192(pi0192),
    .pi0193(pi0193),
    .pi0194(pi0194),
    .pi0195(pi0195),
    .pi0196(pi0196),
    .pi0197(pi0197),
    .pi0198(pi0198),
    .pi0199(pi0199),
    .pi0200(pi0200),
    .pi0201(pi0201),
    .pi0202(pi0202),
    .pi0203(pi0203),
    .pi0204(pi0204),
    .pi0205(pi0205),
    .pi0206(pi0206),
    .pi0207(pi0207),
    .pi0208(pi0208),
    .pi0209(pi0209),
    .pi0210(pi0210),
    .pi0211(pi0211),
    .pi0212(pi0212),
    .pi0213(pi0213),
    .pi0214(pi0214),
    .pi0215(pi0215),
    .pi0216(pi0216),
    .pi0217(pi0217),
    .pi0218(pi0218),
    .pi0219(pi0219),
    .pi0220(pi0220),
    .pi0221(pi0221),
    .pi0222(pi0222),
    .pi0223(pi0223),
    .pi0224(pi0224),
    .pi0225(pi0225),
    .pi0226(pi0226),
    .pi0227(pi0227),
    .pi0228(pi0228),
    .pi0229(pi0229),
    .pi0230(pi0230),
    .pi0231(pi0231),
    .pi0232(pi0232),
    .pi0233(pi0233),
    .pi0234(pi0234),
    .pi0235(pi0235),
    .pi0236(pi0236),
    .pi0237(pi0237),
    .pi0238(pi0238),
    .pi0239(pi0239),
    .pi0240(pi0240),
    .pi0241(pi0241),
    .pi0242(pi0242),
    .pi0243(pi0243),
    .pi0244(pi0244),
    .pi0245(pi0245),
    .pi0246(pi0246),
    .pi0247(pi0247),
    .pi0248(pi0248),
    .pi0249(pi0249),
    .pi0250(pi0250),
    .pi0251(pi0251),
    .pi0252(pi0252),
    .pi0253(pi0253),
    .pi0254(pi0254),
    .pi0255(pi0255),
    .pi0256(pi0256),
    .pi0257(pi0257),
    .pi0258(pi0258),
    .pi0259(pi0259),
    .pi0260(pi0260),
    .pi0261(pi0261),
    .pi0262(pi0262),
    .pi0263(pi0263),
    .pi0264(pi0264),
    .pi0265(pi0265),
    .pi0266(pi0266),
    .pi0267(pi0267),
    .pi0268(pi0268),
    .pi0269(pi0269),
    .pi0270(pi0270),
    .pi0271(pi0271),
    .pi0272(pi0272),
    .pi0273(pi0273),
    .pi0274(pi0274),
    .pi0275(pi0275),
    .pi0276(pi0276),
    .pi0277(pi0277),
    .pi0278(pi0278),
    .pi0279(pi0279),
    .pi0280(pi0280),
    .pi0281(pi0281),
    .pi0282(pi0282),
    .pi0283(pi0283),
    .pi0284(pi0284),
    .pi0285(pi0285),
    .pi0286(pi0286),
    .pi0287(pi0287),
    .pi0288(pi0288),
    .pi0289(pi0289),
    .pi0290(pi0290),
    .pi0291(pi0291),
    .pi0292(pi0292),
    .pi0293(pi0293),
    .pi0294(pi0294),
    .pi0295(pi0295),
    .pi0296(pi0296),
    .pi0297(pi0297),
    .pi0298(pi0298),
    .pi0299(pi0299),
    .pi0300(pi0300),
    .pi0301(pi0301),
    .pi0302(pi0302),
    .pi0303(pi0303),
    .pi0304(pi0304),
    .pi0305(pi0305),
    .pi0306(pi0306),
    .pi0307(pi0307),
    .pi0308(pi0308),
    .pi0309(pi0309),
    .pi0310(pi0310),
    .pi0311(pi0311),
    .pi0312(pi0312),
    .pi0313(pi0313),
    .pi0314(pi0314),
    .pi0315(pi0315),
    .pi0316(pi0316),
    .pi0317(pi0317),
    .pi0318(pi0318),
    .pi0319(pi0319),
    .pi0320(pi0320),
    .pi0321(pi0321),
    .pi0322(pi0322),
    .pi0323(pi0323),
    .pi0324(pi0324),
    .pi0325(pi0325),
    .pi0326(pi0326),
    .pi0327(pi0327),
    .pi0328(pi0328),
    .pi0329(pi0329),
    .pi0330(pi0330),
    .pi0331(pi0331),
    .pi0332(pi0332),
    .pi0333(pi0333),
    .pi0334(pi0334),
    .pi0335(pi0335),
    .pi0336(pi0336),
    .pi0337(pi0337),
    .pi0338(pi0338),
    .pi0339(pi0339),
    .pi0340(pi0340),
    .pi0341(pi0341),
    .pi0342(pi0342),
    .pi0343(pi0343),
    .pi0344(pi0344),
    .pi0345(pi0345),
    .pi0346(pi0346),
    .pi0347(pi0347),
    .pi0348(pi0348),
    .pi0349(pi0349),
    .pi0350(pi0350),
    .pi0351(pi0351),
    .pi0352(pi0352),
    .pi0353(pi0353),
    .pi0354(pi0354),
    .pi0355(pi0355),
    .pi0356(pi0356),
    .pi0357(pi0357),
    .pi0358(pi0358),
    .pi0359(pi0359),
    .pi0360(pi0360),
    .pi0361(pi0361),
    .pi0362(pi0362),
    .pi0363(pi0363),
    .pi0364(pi0364),
    .pi0365(pi0365),
    .pi0366(pi0366),
    .pi0367(pi0367),
    .pi0368(pi0368),
    .pi0369(pi0369),
    .pi0370(pi0370),
    .pi0371(pi0371),
    .pi0372(pi0372),
    .pi0373(pi0373),
    .pi0374(pi0374),
    .pi0375(pi0375),
    .pi0376(pi0376),
    .pi0377(pi0377),
    .pi0378(pi0378),
    .pi0379(pi0379),
    .pi0380(pi0380),
    .pi0381(pi0381),
    .pi0382(pi0382),
    .pi0383(pi0383),
    .pi0384(pi0384),
    .pi0385(pi0385),
    .pi0386(pi0386),
    .pi0387(pi0387),
    .pi0388(pi0388),
    .pi0389(pi0389),
    .pi0390(pi0390),
    .pi0391(pi0391),
    .pi0392(pi0392),
    .pi0393(pi0393),
    .pi0394(pi0394),
    .pi0395(pi0395),
    .pi0396(pi0396),
    .pi0397(pi0397),
    .pi0398(pi0398),
    .pi0399(pi0399),
    .pi0400(pi0400),
    .pi0401(pi0401),
    .pi0402(pi0402),
    .pi0403(pi0403),
    .pi0404(pi0404),
    .pi0405(pi0405),
    .pi0406(pi0406),
    .pi0407(pi0407),
    .pi0408(pi0408),
    .pi0409(pi0409),
    .pi0410(pi0410),
    .pi0411(pi0411),
    .pi0412(pi0412),
    .pi0413(pi0413),
    .pi0414(pi0414),
    .pi0415(pi0415),
    .pi0416(pi0416),
    .pi0417(pi0417),
    .pi0418(pi0418),
    .pi0419(pi0419),
    .pi0420(pi0420),
    .pi0421(pi0421),
    .pi0422(pi0422),
    .pi0423(pi0423),
    .pi0424(pi0424),
    .pi0425(pi0425),
    .pi0426(pi0426),
    .pi0427(pi0427),
    .pi0428(pi0428),
    .pi0429(pi0429),
    .pi0430(pi0430),
    .pi0431(pi0431),
    .pi0432(pi0432),
    .pi0433(pi0433),
    .pi0434(pi0434),
    .pi0435(pi0435),
    .pi0436(pi0436),
    .pi0437(pi0437),
    .pi0438(pi0438),
    .pi0439(pi0439),
    .pi0440(pi0440),
    .pi0441(pi0441),
    .pi0442(pi0442),
    .pi0443(pi0443),
    .pi0444(pi0444),
    .pi0445(pi0445),
    .pi0446(pi0446),
    .pi0447(pi0447),
    .pi0448(pi0448),
    .pi0449(pi0449),
    .pi0450(pi0450),
    .pi0451(pi0451),
    .pi0452(pi0452),
    .pi0453(pi0453),
    .pi0454(pi0454),
    .pi0455(pi0455),
    .pi0456(pi0456),
    .pi0457(pi0457),
    .pi0458(pi0458),
    .pi0459(pi0459),
    .pi0460(pi0460),
    .pi0461(pi0461),
    .pi0462(pi0462),
    .pi0463(pi0463),
    .pi0464(pi0464),
    .pi0465(pi0465),
    .pi0466(pi0466),
    .pi0467(pi0467),
    .pi0468(pi0468),
    .pi0469(pi0469),
    .pi0470(pi0470),
    .pi0471(pi0471),
    .pi0472(pi0472),
    .pi0473(pi0473),
    .pi0474(pi0474),
    .pi0475(pi0475),
    .pi0476(pi0476),
    .pi0477(pi0477),
    .pi0478(pi0478),
    .pi0479(pi0479),
    .pi0480(pi0480),
    .pi0481(pi0481),
    .pi0482(pi0482),
    .pi0483(pi0483),
    .pi0484(pi0484),
    .pi0485(pi0485),
    .pi0486(pi0486),
    .pi0487(pi0487),
    .pi0488(pi0488),
    .pi0489(pi0489),
    .pi0490(pi0490),
    .pi0491(pi0491),
    .pi0492(pi0492),
    .pi0493(pi0493),
    .pi0494(pi0494),
    .pi0495(pi0495),
    .pi0496(pi0496),
    .pi0497(pi0497),
    .pi0498(pi0498),
    .pi0499(pi0499),
    .pi0500(pi0500),
    .pi0501(pi0501),
    .pi0502(pi0502),
    .pi0503(pi0503),
    .pi0504(pi0504),
    .pi0505(pi0505),
    .pi0506(pi0506),
    .pi0507(pi0507),
    .pi0508(pi0508),
    .pi0509(pi0509),
    .pi0510(pi0510),
    .pi0511(pi0511),
    .pi0512(pi0512),
    .pi0513(pi0513),
    .pi0514(pi0514),
    .pi0515(pi0515),
    .pi0516(pi0516),
    .pi0517(pi0517),
    .pi0518(pi0518),
    .pi0519(pi0519),
    .pi0520(pi0520),
    .pi0521(pi0521),
    .pi0522(pi0522),
    .pi0523(pi0523),
    .pi0524(pi0524),
    .pi0525(pi0525),
    .pi0526(pi0526),
    .pi0527(pi0527),
    .pi0528(pi0528),
    .pi0529(pi0529),
    .pi0530(pi0530),
    .pi0531(pi0531),
    .pi0532(pi0532),
    .pi0533(pi0533),
    .pi0534(pi0534),
    .pi0535(pi0535),
    .pi0536(pi0536),
    .pi0537(pi0537),
    .pi0538(pi0538),
    .pi0539(pi0539),
    .pi0540(pi0540),
    .pi0541(pi0541),
    .pi0542(pi0542),
    .pi0543(pi0543),
    .pi0544(pi0544),
    .pi0545(pi0545),
    .pi0546(pi0546),
    .pi0547(pi0547),
    .pi0548(pi0548),
    .pi0549(pi0549),
    .pi0550(pi0550),
    .pi0551(pi0551),
    .pi0552(pi0552),
    .pi0553(pi0553),
    .pi0554(pi0554),
    .pi0555(pi0555),
    .pi0556(pi0556),
    .pi0557(pi0557),
    .pi0558(pi0558),
    .pi0559(pi0559),
    .pi0560(pi0560),
    .pi0561(pi0561),
    .pi0562(pi0562),
    .pi0563(pi0563),
    .pi0564(pi0564),
    .pi0565(pi0565),
    .pi0566(pi0566),
    .pi0567(pi0567),
    .pi0568(pi0568),
    .pi0569(pi0569),
    .pi0570(pi0570),
    .pi0571(pi0571),
    .pi0572(pi0572),
    .pi0573(pi0573),
    .pi0574(pi0574),
    .pi0575(pi0575),
    .pi0576(pi0576),
    .pi0577(pi0577),
    .pi0578(pi0578),
    .pi0579(pi0579),
    .pi0580(pi0580),
    .pi0581(pi0581),
    .pi0582(pi0582),
    .pi0583(pi0583),
    .pi0584(pi0584),
    .pi0585(pi0585),
    .pi0586(pi0586),
    .pi0587(pi0587),
    .pi0588(pi0588),
    .pi0589(pi0589),
    .pi0590(pi0590),
    .pi0591(pi0591),
    .pi0592(pi0592),
    .pi0593(pi0593),
    .pi0594(pi0594),
    .pi0595(pi0595),
    .pi0596(pi0596),
    .pi0597(pi0597),
    .pi0598(pi0598),
    .pi0599(pi0599),
    .pi0600(pi0600),
    .pi0601(pi0601),
    .pi0602(pi0602),
    .pi0603(pi0603),
    .pi0604(pi0604),
    .pi0605(pi0605),
    .pi0606(pi0606),
    .pi0607(pi0607),
    .pi0608(pi0608),
    .pi0609(pi0609),
    .pi0610(pi0610),
    .pi0611(pi0611),
    .pi0612(pi0612),
    .pi0613(pi0613),
    .pi0614(pi0614),
    .pi0615(pi0615),
    .pi0616(pi0616),
    .pi0617(pi0617),
    .pi0618(pi0618),
    .pi0619(pi0619),
    .pi0620(pi0620),
    .pi0621(pi0621),
    .pi0622(pi0622),
    .pi0623(pi0623),
    .pi0624(pi0624),
    .pi0625(pi0625),
    .pi0626(pi0626),
    .pi0627(pi0627),
    .pi0628(pi0628),
    .pi0629(pi0629),
    .pi0630(pi0630),
    .pi0631(pi0631),
    .pi0632(pi0632),
    .pi0633(pi0633),
    .pi0634(pi0634),
    .pi0635(pi0635),
    .pi0636(pi0636),
    .pi0637(pi0637),
    .pi0638(pi0638),
    .pi0639(pi0639),
    .pi0640(pi0640),
    .pi0641(pi0641),
    .pi0642(pi0642),
    .pi0643(pi0643),
    .pi0644(pi0644),
    .pi0645(pi0645),
    .pi0646(pi0646),
    .pi0647(pi0647),
    .pi0648(pi0648),
    .pi0649(pi0649),
    .pi0650(pi0650),
    .pi0651(pi0651),
    .pi0652(pi0652),
    .pi0653(pi0653),
    .pi0654(pi0654),
    .pi0655(pi0655),
    .pi0656(pi0656),
    .pi0657(pi0657),
    .pi0658(pi0658),
    .pi0659(pi0659),
    .pi0660(pi0660),
    .pi0661(pi0661),
    .pi0662(pi0662),
    .pi0663(pi0663),
    .pi0664(pi0664),
    .pi0665(pi0665),
    .pi0666(pi0666),
    .pi0667(pi0667),
    .pi0668(pi0668),
    .pi0669(pi0669),
    .pi0670(pi0670),
    .pi0671(pi0671),
    .pi0672(pi0672),
    .pi0673(pi0673),
    .pi0674(pi0674),
    .pi0675(pi0675),
    .pi0676(pi0676),
    .pi0677(pi0677),
    .pi0678(pi0678),
    .pi0679(pi0679),
    .pi0680(pi0680),
    .pi0681(pi0681),
    .pi0682(pi0682),
    .pi0683(pi0683),
    .pi0684(pi0684),
    .pi0685(pi0685),
    .pi0686(pi0686),
    .pi0687(pi0687),
    .pi0688(pi0688),
    .pi0689(pi0689),
    .pi0690(pi0690),
    .pi0691(pi0691),
    .pi0692(pi0692),
    .pi0693(pi0693),
    .pi0694(pi0694),
    .pi0695(pi0695),
    .pi0696(pi0696),
    .pi0697(pi0697),
    .pi0698(pi0698),
    .pi0699(pi0699),
    .pi0700(pi0700),
    .pi0701(pi0701),
    .pi0702(pi0702),
    .pi0703(pi0703),
    .pi0704(pi0704),
    .pi0705(pi0705),
    .pi0706(pi0706),
    .pi0707(pi0707),
    .pi0708(pi0708),
    .pi0709(pi0709),
    .pi0710(pi0710),
    .pi0711(pi0711),
    .pi0712(pi0712),
    .pi0713(pi0713),
    .pi0714(pi0714),
    .pi0715(pi0715),
    .pi0716(pi0716),
    .pi0717(pi0717),
    .pi0718(pi0718),
    .pi0719(pi0719),
    .pi0720(pi0720),
    .pi0721(pi0721),
    .pi0722(pi0722),
    .pi0723(pi0723),
    .pi0724(pi0724),
    .pi0725(pi0725),
    .pi0726(pi0726),
    .pi0727(pi0727),
    .pi0728(pi0728),
    .pi0729(pi0729),
    .pi0730(pi0730),
    .pi0731(pi0731),
    .pi0732(pi0732),
    .pi0733(pi0733),
    .pi0734(pi0734),
    .pi0735(pi0735),
    .pi0736(pi0736),
    .pi0737(pi0737),
    .pi0738(pi0738),
    .pi0739(pi0739),
    .pi0740(pi0740),
    .pi0741(pi0741),
    .pi0742(pi0742),
    .pi0743(pi0743),
    .pi0744(pi0744),
    .pi0745(pi0745),
    .pi0746(pi0746),
    .pi0747(pi0747),
    .pi0748(pi0748),
    .pi0749(pi0749),
    .pi0750(pi0750),
    .pi0751(pi0751),
    .pi0752(pi0752),
    .pi0753(pi0753),
    .pi0754(pi0754),
    .pi0755(pi0755),
    .pi0756(pi0756),
    .pi0757(pi0757),
    .pi0758(pi0758),
    .pi0759(pi0759),
    .pi0760(pi0760),
    .pi0761(pi0761),
    .pi0762(pi0762),
    .pi0763(pi0763),
    .pi0764(pi0764),
    .pi0765(pi0765),
    .pi0766(pi0766),
    .pi0767(pi0767),
    .pi0768(pi0768),
    .pi0769(pi0769),
    .pi0770(pi0770),
    .pi0771(pi0771),
    .pi0772(pi0772),
    .pi0773(pi0773),
    .pi0774(pi0774),
    .pi0775(pi0775),
    .pi0776(pi0776),
    .pi0777(pi0777),
    .pi0778(pi0778),
    .pi0779(pi0779),
    .pi0780(pi0780),
    .pi0781(pi0781),
    .pi0782(pi0782),
    .pi0783(pi0783),
    .pi0784(pi0784),
    .pi0785(pi0785),
    .pi0786(pi0786),
    .pi0787(pi0787),
    .pi0788(pi0788),
    .pi0789(pi0789),
    .pi0790(pi0790),
    .pi0791(pi0791),
    .pi0792(pi0792),
    .pi0793(pi0793),
    .pi0794(pi0794),
    .pi0795(pi0795),
    .pi0796(pi0796),
    .pi0797(pi0797),
    .pi0798(pi0798),
    .pi0799(pi0799),
    .pi0800(pi0800),
    .pi0801(pi0801),
    .pi0802(pi0802),
    .pi0803(pi0803),
    .pi0804(pi0804),
    .pi0805(pi0805),
    .pi0806(pi0806),
    .pi0807(pi0807),
    .pi0808(pi0808),
    .pi0809(pi0809),
    .pi0810(pi0810),
    .pi0811(pi0811),
    .pi0812(pi0812),
    .pi0813(pi0813),
    .pi0814(pi0814),
    .pi0815(pi0815),
    .pi0816(pi0816),
    .pi0817(pi0817),
    .pi0818(pi0818),
    .pi0819(pi0819),
    .pi0820(pi0820),
    .pi0821(pi0821),
    .pi0822(pi0822),
    .pi0823(pi0823),
    .pi0824(pi0824),
    .pi0825(pi0825),
    .pi0826(pi0826),
    .pi0827(pi0827),
    .pi0828(pi0828),
    .pi0829(pi0829),
    .pi0830(pi0830),
    .pi0831(pi0831),
    .pi0832(pi0832),
    .pi0833(pi0833),
    .pi0834(pi0834),
    .pi0835(pi0835),
    .pi0836(pi0836),
    .pi0837(pi0837),
    .pi0838(pi0838),
    .pi0839(pi0839),
    .pi0840(pi0840),
    .pi0841(pi0841),
    .pi0842(pi0842),
    .pi0843(pi0843),
    .pi0844(pi0844),
    .pi0845(pi0845),
    .pi0846(pi0846),
    .pi0847(pi0847),
    .pi0848(pi0848),
    .pi0849(pi0849),
    .pi0850(pi0850),
    .pi0851(pi0851),
    .pi0852(pi0852),
    .pi0853(pi0853),
    .pi0854(pi0854),
    .pi0855(pi0855),
    .pi0856(pi0856),
    .pi0857(pi0857),
    .pi0858(pi0858),
    .pi0859(pi0859),
    .pi0860(pi0860),
    .pi0861(pi0861),
    .pi0862(pi0862),
    .pi0863(pi0863),
    .pi0864(pi0864),
    .pi0865(pi0865),
    .pi0866(pi0866),
    .pi0867(pi0867),
    .pi0868(pi0868),
    .pi0869(pi0869),
    .pi0870(pi0870),
    .pi0871(pi0871),
    .pi0872(pi0872),
    .pi0873(pi0873),
    .pi0874(pi0874),
    .pi0875(pi0875),
    .pi0876(pi0876),
    .pi0877(pi0877),
    .pi0878(pi0878),
    .pi0879(pi0879),
    .pi0880(pi0880),
    .pi0881(pi0881),
    .pi0882(pi0882),
    .pi0883(pi0883),
    .pi0884(pi0884),
    .pi0885(pi0885),
    .pi0886(pi0886),
    .pi0887(pi0887),
    .pi0888(pi0888),
    .pi0889(pi0889),
    .pi0890(pi0890),
    .pi0891(pi0891),
    .pi0892(pi0892),
    .pi0893(pi0893),
    .pi0894(pi0894),
    .pi0895(pi0895),
    .pi0896(pi0896),
    .pi0897(pi0897),
    .pi0898(pi0898),
    .pi0899(pi0899),
    .pi0900(pi0900),
    .pi0901(pi0901),
    .pi0902(pi0902),
    .pi0903(pi0903),
    .pi0904(pi0904),
    .pi0905(pi0905),
    .pi0906(pi0906),
    .pi0907(pi0907),
    .pi0908(pi0908),
    .pi0909(pi0909),
    .pi0910(pi0910),
    .pi0911(pi0911),
    .pi0912(pi0912),
    .pi0913(pi0913),
    .pi0914(pi0914),
    .pi0915(pi0915),
    .pi0916(pi0916),
    .pi0917(pi0917),
    .pi0918(pi0918),
    .pi0919(pi0919),
    .pi0920(pi0920),
    .pi0921(pi0921),
    .pi0922(pi0922),
    .pi0923(pi0923),
    .pi0924(pi0924),
    .pi0925(pi0925),
    .pi0926(pi0926),
    .pi0927(pi0927),
    .pi0928(pi0928),
    .pi0929(pi0929),
    .pi0930(pi0930),
    .pi0931(pi0931),
    .pi0932(pi0932),
    .pi0933(pi0933),
    .pi0934(pi0934),
    .pi0935(pi0935),
    .pi0936(pi0936),
    .pi0937(pi0937),
    .pi0938(pi0938),
    .pi0939(pi0939),
    .pi0940(pi0940),
    .pi0941(pi0941),
    .pi0942(pi0942),
    .pi0943(pi0943),
    .pi0944(pi0944),
    .pi0945(pi0945),
    .pi0946(pi0946),
    .pi0947(pi0947),
    .pi0948(pi0948),
    .pi0949(pi0949),
    .pi0950(pi0950),
    .pi0951(pi0951),
    .pi0952(pi0952),
    .pi0953(pi0953),
    .pi0954(pi0954),
    .pi0955(pi0955),
    .pi0956(pi0956),
    .pi0957(pi0957),
    .pi0958(pi0958),
    .pi0959(pi0959),
    .pi0960(pi0960),
    .pi0961(pi0961),
    .pi0962(pi0962),
    .pi0963(pi0963),
    .pi0964(pi0964),
    .pi0965(pi0965),
    .pi0966(pi0966),
    .pi0967(pi0967),
    .pi0968(pi0968),
    .pi0969(pi0969),
    .pi0970(pi0970),
    .pi0971(pi0971),
    .pi0972(pi0972),
    .pi0973(pi0973),
    .pi0974(pi0974),
    .pi0975(pi0975),
    .pi0976(pi0976),
    .pi0977(pi0977),
    .pi0978(pi0978),
    .pi0979(pi0979),
    .pi0980(pi0980),
    .pi0981(pi0981),
    .pi0982(pi0982),
    .pi0983(pi0983),
    .pi0984(pi0984),
    .pi0985(pi0985),
    .pi0986(pi0986),
    .pi0987(pi0987),
    .pi0988(pi0988),
    .pi0989(pi0989),
    .pi0990(pi0990),
    .pi0991(pi0991),
    .pi0992(pi0992),
    .pi0993(pi0993),
    .pi0994(pi0994),
    .pi0995(pi0995),
    .pi0996(pi0996),
    .pi0997(pi0997),
    .pi0998(pi0998),
    .pi0999(pi0999),
    .pi1000(pi1000),
    .pi1001(pi1001),
    .pi1002(pi1002),
    .pi1003(pi1003),
    .pi1004(pi1004),
    .pi1005(pi1005),
    .pi1006(pi1006),
    .pi1007(pi1007),
    .pi1008(pi1008),
    .pi1009(pi1009),
    .pi1010(pi1010),
    .pi1011(pi1011),
    .pi1012(pi1012),
    .pi1013(pi1013),
    .pi1014(pi1014),
    .pi1015(pi1015),
    .pi1016(pi1016),
    .pi1017(pi1017),
    .pi1018(pi1018),
    .pi1019(pi1019),
    .pi1020(pi1020),
    .pi1021(pi1021),
    .pi1022(pi1022),
    .pi1023(pi1023),
    .pi1024(pi1024),
    .pi1025(pi1025),
    .pi1026(pi1026),
    .pi1027(pi1027),
    .pi1028(pi1028),
    .pi1029(pi1029),
    .pi1030(pi1030),
    .pi1031(pi1031),
    .pi1032(pi1032),
    .pi1033(pi1033),
    .pi1034(pi1034),
    .pi1035(pi1035),
    .pi1036(pi1036),
    .pi1037(pi1037),
    .pi1038(pi1038),
    .pi1039(pi1039),
    .pi1040(pi1040),
    .pi1041(pi1041),
    .pi1042(pi1042),
    .pi1043(pi1043),
    .pi1044(pi1044),
    .pi1045(pi1045),
    .pi1046(pi1046),
    .pi1047(pi1047),
    .pi1048(pi1048),
    .pi1049(pi1049),
    .pi1050(pi1050),
    .pi1051(pi1051),
    .pi1052(pi1052),
    .pi1053(pi1053),
    .pi1054(pi1054),
    .pi1055(pi1055),
    .pi1056(pi1056),
    .pi1057(pi1057),
    .pi1058(pi1058),
    .pi1059(pi1059),
    .pi1060(pi1060),
    .pi1061(pi1061),
    .pi1062(pi1062),
    .pi1063(pi1063),
    .pi1064(pi1064),
    .pi1065(pi1065),
    .pi1066(pi1066),
    .pi1067(pi1067),
    .pi1068(pi1068),
    .pi1069(pi1069),
    .pi1070(pi1070),
    .pi1071(pi1071),
    .pi1072(pi1072),
    .pi1073(pi1073),
    .pi1074(pi1074),
    .pi1075(pi1075),
    .pi1076(pi1076),
    .pi1077(pi1077),
    .pi1078(pi1078),
    .pi1079(pi1079),
    .pi1080(pi1080),
    .pi1081(pi1081),
    .pi1082(pi1082),
    .pi1083(pi1083),
    .pi1084(pi1084),
    .pi1085(pi1085),
    .pi1086(pi1086),
    .pi1087(pi1087),
    .pi1088(pi1088),
    .pi1089(pi1089),
    .pi1090(pi1090),
    .pi1091(pi1091),
    .pi1092(pi1092),
    .pi1093(pi1093),
    .pi1094(pi1094),
    .pi1095(pi1095),
    .pi1096(pi1096),
    .pi1097(pi1097),
    .pi1098(pi1098),
    .pi1099(pi1099),
    .pi1100(pi1100),
    .pi1101(pi1101),
    .pi1102(pi1102),
    .pi1103(pi1103),
    .pi1104(pi1104),
    .pi1105(pi1105),
    .pi1106(pi1106),
    .pi1107(pi1107),
    .pi1108(pi1108),
    .pi1109(pi1109),
    .pi1110(pi1110),
    .pi1111(pi1111),
    .pi1112(pi1112),
    .pi1113(pi1113),
    .pi1114(pi1114),
    .pi1115(pi1115),
    .pi1116(pi1116),
    .pi1117(pi1117),
    .pi1118(pi1118),
    .pi1119(pi1119),
    .pi1120(pi1120),
    .pi1121(pi1121),
    .pi1122(pi1122),
    .pi1123(pi1123),
    .pi1124(pi1124),
    .pi1125(pi1125),
    .pi1126(pi1126),
    .pi1127(pi1127),
    .pi1128(pi1128),
    .pi1129(pi1129),
    .pi1130(pi1130),
    .pi1131(pi1131),
    .pi1132(pi1132),
    .pi1133(pi1133),
    .pi1134(pi1134),
    .pi1135(pi1135),
    .pi1136(pi1136),
    .pi1137(pi1137),
    .pi1138(pi1138),
    .pi1139(pi1139),
    .pi1140(pi1140),
    .pi1141(pi1141),
    .pi1142(pi1142),
    .pi1143(pi1143),
    .pi1144(pi1144),
    .pi1145(pi1145),
    .pi1146(pi1146),
    .pi1147(pi1147),
    .pi1148(pi1148),
    .pi1149(pi1149),
    .pi1150(pi1150),
    .pi1151(pi1151),
    .pi1152(pi1152),
    .pi1153(pi1153),
    .pi1154(pi1154),
    .pi1155(pi1155),
    .pi1156(pi1156),
    .pi1157(pi1157),
    .pi1158(pi1158),
    .pi1159(pi1159),
    .pi1160(pi1160),
    .pi1161(pi1161),
    .pi1162(pi1162),
    .pi1163(pi1163),
    .pi1164(pi1164),
    .pi1165(pi1165),
    .pi1166(pi1166),
    .pi1167(pi1167),
    .pi1168(pi1168),
    .pi1169(pi1169),
    .pi1170(pi1170),
    .pi1171(pi1171),
    .pi1172(pi1172),
    .pi1173(pi1173),
    .pi1174(pi1174),
    .pi1175(pi1175),
    .pi1176(pi1176),
    .pi1177(pi1177),
    .pi1178(pi1178),
    .pi1179(pi1179),
    .pi1180(pi1180),
    .pi1181(pi1181),
    .pi1182(pi1182),
    .pi1183(pi1183),
    .pi1184(pi1184),
    .pi1185(pi1185),
    .pi1186(pi1186),
    .pi1187(pi1187),
    .pi1188(pi1188),
    .pi1189(pi1189),
    .pi1190(pi1190),
    .pi1191(pi1191),
    .pi1192(pi1192),
    .pi1193(pi1193),
    .pi1194(pi1194),
    .pi1195(pi1195),
    .pi1196(pi1196),
    .pi1197(pi1197),
    .pi1198(pi1198),
    .pi1199(pi1199),
    .pi1200(pi1200),
    .pi1201(pi1201),
    .pi1202(pi1202),
    .pi1203(pi1203),
    .po0000(po0000),
    .po0001(po0001),
    .po0002(po0002),
    .po0003(po0003),
    .po0004(po0004),
    .po0005(po0005),
    .po0006(po0006),
    .po0007(po0007),
    .po0008(po0008),
    .po0009(po0009),
    .po0010(po0010),
    .po0011(po0011),
    .po0012(po0012),
    .po0013(po0013),
    .po0014(po0014),
    .po0015(po0015),
    .po0016(po0016),
    .po0017(po0017),
    .po0018(po0018),
    .po0019(po0019),
    .po0020(po0020),
    .po0021(po0021),
    .po0022(po0022),
    .po0023(po0023),
    .po0024(po0024),
    .po0025(po0025),
    .po0026(po0026),
    .po0027(po0027),
    .po0028(po0028),
    .po0029(po0029),
    .po0030(po0030),
    .po0031(po0031),
    .po0032(po0032),
    .po0033(po0033),
    .po0034(po0034),
    .po0035(po0035),
    .po0036(po0036),
    .po0037(po0037),
    .po0038(po0038),
    .po0039(po0039),
    .po0040(po0040),
    .po0041(po0041),
    .po0042(po0042),
    .po0043(po0043),
    .po0044(po0044),
    .po0045(po0045),
    .po0046(po0046),
    .po0047(po0047),
    .po0048(po0048),
    .po0049(po0049),
    .po0050(po0050),
    .po0051(po0051),
    .po0052(po0052),
    .po0053(po0053),
    .po0054(po0054),
    .po0055(po0055),
    .po0056(po0056),
    .po0057(po0057),
    .po0058(po0058),
    .po0059(po0059),
    .po0060(po0060),
    .po0061(po0061),
    .po0062(po0062),
    .po0063(po0063),
    .po0064(po0064),
    .po0065(po0065),
    .po0066(po0066),
    .po0067(po0067),
    .po0068(po0068),
    .po0069(po0069),
    .po0070(po0070),
    .po0071(po0071),
    .po0072(po0072),
    .po0073(po0073),
    .po0074(po0074),
    .po0075(po0075),
    .po0076(po0076),
    .po0077(po0077),
    .po0078(po0078),
    .po0079(po0079),
    .po0080(po0080),
    .po0081(po0081),
    .po0082(po0082),
    .po0083(po0083),
    .po0084(po0084),
    .po0085(po0085),
    .po0086(po0086),
    .po0087(po0087),
    .po0088(po0088),
    .po0089(po0089),
    .po0090(po0090),
    .po0091(po0091),
    .po0092(po0092),
    .po0093(po0093),
    .po0094(po0094),
    .po0095(po0095),
    .po0096(po0096),
    .po0097(po0097),
    .po0098(po0098),
    .po0099(po0099),
    .po0100(po0100),
    .po0101(po0101),
    .po0102(po0102),
    .po0103(po0103),
    .po0104(po0104),
    .po0105(po0105),
    .po0106(po0106),
    .po0107(po0107),
    .po0108(po0108),
    .po0109(po0109),
    .po0110(po0110),
    .po0111(po0111),
    .po0112(po0112),
    .po0113(po0113),
    .po0114(po0114),
    .po0115(po0115),
    .po0116(po0116),
    .po0117(po0117),
    .po0118(po0118),
    .po0119(po0119),
    .po0120(po0120),
    .po0121(po0121),
    .po0122(po0122),
    .po0123(po0123),
    .po0124(po0124),
    .po0125(po0125),
    .po0126(po0126),
    .po0127(po0127),
    .po0128(po0128),
    .po0129(po0129),
    .po0130(po0130),
    .po0131(po0131),
    .po0132(po0132),
    .po0133(po0133),
    .po0134(po0134),
    .po0135(po0135),
    .po0136(po0136),
    .po0137(po0137),
    .po0138(po0138),
    .po0139(po0139),
    .po0140(po0140),
    .po0141(po0141),
    .po0142(po0142),
    .po0143(po0143),
    .po0144(po0144),
    .po0145(po0145),
    .po0146(po0146),
    .po0147(po0147),
    .po0148(po0148),
    .po0149(po0149),
    .po0150(po0150),
    .po0151(po0151),
    .po0152(po0152),
    .po0153(po0153),
    .po0154(po0154),
    .po0155(po0155),
    .po0156(po0156),
    .po0157(po0157),
    .po0158(po0158),
    .po0159(po0159),
    .po0160(po0160),
    .po0161(po0161),
    .po0162(po0162),
    .po0163(po0163),
    .po0164(po0164),
    .po0165(po0165),
    .po0166(po0166),
    .po0167(po0167),
    .po0168(po0168),
    .po0169(po0169),
    .po0170(po0170),
    .po0171(po0171),
    .po0172(po0172),
    .po0173(po0173),
    .po0174(po0174),
    .po0175(po0175),
    .po0176(po0176),
    .po0177(po0177),
    .po0178(po0178),
    .po0179(po0179),
    .po0180(po0180),
    .po0181(po0181),
    .po0182(po0182),
    .po0183(po0183),
    .po0184(po0184),
    .po0185(po0185),
    .po0186(po0186),
    .po0187(po0187),
    .po0188(po0188),
    .po0189(po0189),
    .po0190(po0190),
    .po0191(po0191),
    .po0192(po0192),
    .po0193(po0193),
    .po0194(po0194),
    .po0195(po0195),
    .po0196(po0196),
    .po0197(po0197),
    .po0198(po0198),
    .po0199(po0199),
    .po0200(po0200),
    .po0201(po0201),
    .po0202(po0202),
    .po0203(po0203),
    .po0204(po0204),
    .po0205(po0205),
    .po0206(po0206),
    .po0207(po0207),
    .po0208(po0208),
    .po0209(po0209),
    .po0210(po0210),
    .po0211(po0211),
    .po0212(po0212),
    .po0213(po0213),
    .po0214(po0214),
    .po0215(po0215),
    .po0216(po0216),
    .po0217(po0217),
    .po0218(po0218),
    .po0219(po0219),
    .po0220(po0220),
    .po0221(po0221),
    .po0222(po0222),
    .po0223(po0223),
    .po0224(po0224),
    .po0225(po0225),
    .po0226(po0226),
    .po0227(po0227),
    .po0228(po0228),
    .po0229(po0229),
    .po0230(po0230),
    .po0231(po0231),
    .po0232(po0232),
    .po0233(po0233),
    .po0234(po0234),
    .po0235(po0235),
    .po0236(po0236),
    .po0237(po0237),
    .po0238(po0238),
    .po0239(po0239),
    .po0240(po0240),
    .po0241(po0241),
    .po0242(po0242),
    .po0243(po0243),
    .po0244(po0244),
    .po0245(po0245),
    .po0246(po0246),
    .po0247(po0247),
    .po0248(po0248),
    .po0249(po0249),
    .po0250(po0250),
    .po0251(po0251),
    .po0252(po0252),
    .po0253(po0253),
    .po0254(po0254),
    .po0255(po0255),
    .po0256(po0256),
    .po0257(po0257),
    .po0258(po0258),
    .po0259(po0259),
    .po0260(po0260),
    .po0261(po0261),
    .po0262(po0262),
    .po0263(po0263),
    .po0264(po0264),
    .po0265(po0265),
    .po0266(po0266),
    .po0267(po0267),
    .po0268(po0268),
    .po0269(po0269),
    .po0270(po0270),
    .po0271(po0271),
    .po0272(po0272),
    .po0273(po0273),
    .po0274(po0274),
    .po0275(po0275),
    .po0276(po0276),
    .po0277(po0277),
    .po0278(po0278),
    .po0279(po0279),
    .po0280(po0280),
    .po0281(po0281),
    .po0282(po0282),
    .po0283(po0283),
    .po0284(po0284),
    .po0285(po0285),
    .po0286(po0286),
    .po0287(po0287),
    .po0288(po0288),
    .po0289(po0289),
    .po0290(po0290),
    .po0291(po0291),
    .po0292(po0292),
    .po0293(po0293),
    .po0294(po0294),
    .po0295(po0295),
    .po0296(po0296),
    .po0297(po0297),
    .po0298(po0298),
    .po0299(po0299),
    .po0300(po0300),
    .po0301(po0301),
    .po0302(po0302),
    .po0303(po0303),
    .po0304(po0304),
    .po0305(po0305),
    .po0306(po0306),
    .po0307(po0307),
    .po0308(po0308),
    .po0309(po0309),
    .po0310(po0310),
    .po0311(po0311),
    .po0312(po0312),
    .po0313(po0313),
    .po0314(po0314),
    .po0315(po0315),
    .po0316(po0316),
    .po0317(po0317),
    .po0318(po0318),
    .po0319(po0319),
    .po0320(po0320),
    .po0321(po0321),
    .po0322(po0322),
    .po0323(po0323),
    .po0324(po0324),
    .po0325(po0325),
    .po0326(po0326),
    .po0327(po0327),
    .po0328(po0328),
    .po0329(po0329),
    .po0330(po0330),
    .po0331(po0331),
    .po0332(po0332),
    .po0333(po0333),
    .po0334(po0334),
    .po0335(po0335),
    .po0336(po0336),
    .po0337(po0337),
    .po0338(po0338),
    .po0339(po0339),
    .po0340(po0340),
    .po0341(po0341),
    .po0342(po0342),
    .po0343(po0343),
    .po0344(po0344),
    .po0345(po0345),
    .po0346(po0346),
    .po0347(po0347),
    .po0348(po0348),
    .po0349(po0349),
    .po0350(po0350),
    .po0351(po0351),
    .po0352(po0352),
    .po0353(po0353),
    .po0354(po0354),
    .po0355(po0355),
    .po0356(po0356),
    .po0357(po0357),
    .po0358(po0358),
    .po0359(po0359),
    .po0360(po0360),
    .po0361(po0361),
    .po0362(po0362),
    .po0363(po0363),
    .po0364(po0364),
    .po0365(po0365),
    .po0366(po0366),
    .po0367(po0367),
    .po0368(po0368),
    .po0369(po0369),
    .po0370(po0370),
    .po0371(po0371),
    .po0372(po0372),
    .po0373(po0373),
    .po0374(po0374),
    .po0375(po0375),
    .po0376(po0376),
    .po0377(po0377),
    .po0378(po0378),
    .po0379(po0379),
    .po0380(po0380),
    .po0381(po0381),
    .po0382(po0382),
    .po0383(po0383),
    .po0384(po0384),
    .po0385(po0385),
    .po0386(po0386),
    .po0387(po0387),
    .po0388(po0388),
    .po0389(po0389),
    .po0390(po0390),
    .po0391(po0391),
    .po0392(po0392),
    .po0393(po0393),
    .po0394(po0394),
    .po0395(po0395),
    .po0396(po0396),
    .po0397(po0397),
    .po0398(po0398),
    .po0399(po0399),
    .po0400(po0400),
    .po0401(po0401),
    .po0402(po0402),
    .po0403(po0403),
    .po0404(po0404),
    .po0405(po0405),
    .po0406(po0406),
    .po0407(po0407),
    .po0408(po0408),
    .po0409(po0409),
    .po0410(po0410),
    .po0411(po0411),
    .po0412(po0412),
    .po0413(po0413),
    .po0414(po0414),
    .po0415(po0415),
    .po0416(po0416),
    .po0417(po0417),
    .po0418(po0418),
    .po0419(po0419),
    .po0420(po0420),
    .po0421(po0421),
    .po0422(po0422),
    .po0423(po0423),
    .po0424(po0424),
    .po0425(po0425),
    .po0426(po0426),
    .po0427(po0427),
    .po0428(po0428),
    .po0429(po0429),
    .po0430(po0430),
    .po0431(po0431),
    .po0432(po0432),
    .po0433(po0433),
    .po0434(po0434),
    .po0435(po0435),
    .po0436(po0436),
    .po0437(po0437),
    .po0438(po0438),
    .po0439(po0439),
    .po0440(po0440),
    .po0441(po0441),
    .po0442(po0442),
    .po0443(po0443),
    .po0444(po0444),
    .po0445(po0445),
    .po0446(po0446),
    .po0447(po0447),
    .po0448(po0448),
    .po0449(po0449),
    .po0450(po0450),
    .po0451(po0451),
    .po0452(po0452),
    .po0453(po0453),
    .po0454(po0454),
    .po0455(po0455),
    .po0456(po0456),
    .po0457(po0457),
    .po0458(po0458),
    .po0459(po0459),
    .po0460(po0460),
    .po0461(po0461),
    .po0462(po0462),
    .po0463(po0463),
    .po0464(po0464),
    .po0465(po0465),
    .po0466(po0466),
    .po0467(po0467),
    .po0468(po0468),
    .po0469(po0469),
    .po0470(po0470),
    .po0471(po0471),
    .po0472(po0472),
    .po0473(po0473),
    .po0474(po0474),
    .po0475(po0475),
    .po0476(po0476),
    .po0477(po0477),
    .po0478(po0478),
    .po0479(po0479),
    .po0480(po0480),
    .po0481(po0481),
    .po0482(po0482),
    .po0483(po0483),
    .po0484(po0484),
    .po0485(po0485),
    .po0486(po0486),
    .po0487(po0487),
    .po0488(po0488),
    .po0489(po0489),
    .po0490(po0490),
    .po0491(po0491),
    .po0492(po0492),
    .po0493(po0493),
    .po0494(po0494),
    .po0495(po0495),
    .po0496(po0496),
    .po0497(po0497),
    .po0498(po0498),
    .po0499(po0499),
    .po0500(po0500),
    .po0501(po0501),
    .po0502(po0502),
    .po0503(po0503),
    .po0504(po0504),
    .po0505(po0505),
    .po0506(po0506),
    .po0507(po0507),
    .po0508(po0508),
    .po0509(po0509),
    .po0510(po0510),
    .po0511(po0511),
    .po0512(po0512),
    .po0513(po0513),
    .po0514(po0514),
    .po0515(po0515),
    .po0516(po0516),
    .po0517(po0517),
    .po0518(po0518),
    .po0519(po0519),
    .po0520(po0520),
    .po0521(po0521),
    .po0522(po0522),
    .po0523(po0523),
    .po0524(po0524),
    .po0525(po0525),
    .po0526(po0526),
    .po0527(po0527),
    .po0528(po0528),
    .po0529(po0529),
    .po0530(po0530),
    .po0531(po0531),
    .po0532(po0532),
    .po0533(po0533),
    .po0534(po0534),
    .po0535(po0535),
    .po0536(po0536),
    .po0537(po0537),
    .po0538(po0538),
    .po0539(po0539),
    .po0540(po0540),
    .po0541(po0541),
    .po0542(po0542),
    .po0543(po0543),
    .po0544(po0544),
    .po0545(po0545),
    .po0546(po0546),
    .po0547(po0547),
    .po0548(po0548),
    .po0549(po0549),
    .po0550(po0550),
    .po0551(po0551),
    .po0552(po0552),
    .po0553(po0553),
    .po0554(po0554),
    .po0555(po0555),
    .po0556(po0556),
    .po0557(po0557),
    .po0558(po0558),
    .po0559(po0559),
    .po0560(po0560),
    .po0561(po0561),
    .po0562(po0562),
    .po0563(po0563),
    .po0564(po0564),
    .po0565(po0565),
    .po0566(po0566),
    .po0567(po0567),
    .po0568(po0568),
    .po0569(po0569),
    .po0570(po0570),
    .po0571(po0571),
    .po0572(po0572),
    .po0573(po0573),
    .po0574(po0574),
    .po0575(po0575),
    .po0576(po0576),
    .po0577(po0577),
    .po0578(po0578),
    .po0579(po0579),
    .po0580(po0580),
    .po0581(po0581),
    .po0582(po0582),
    .po0583(po0583),
    .po0584(po0584),
    .po0585(po0585),
    .po0586(po0586),
    .po0587(po0587),
    .po0588(po0588),
    .po0589(po0589),
    .po0590(po0590),
    .po0591(po0591),
    .po0592(po0592),
    .po0593(po0593),
    .po0594(po0594),
    .po0595(po0595),
    .po0596(po0596),
    .po0597(po0597),
    .po0598(po0598),
    .po0599(po0599),
    .po0600(po0600),
    .po0601(po0601),
    .po0602(po0602),
    .po0603(po0603),
    .po0604(po0604),
    .po0605(po0605),
    .po0606(po0606),
    .po0607(po0607),
    .po0608(po0608),
    .po0609(po0609),
    .po0610(po0610),
    .po0611(po0611),
    .po0612(po0612),
    .po0613(po0613),
    .po0614(po0614),
    .po0615(po0615),
    .po0616(po0616),
    .po0617(po0617),
    .po0618(po0618),
    .po0619(po0619),
    .po0620(po0620),
    .po0621(po0621),
    .po0622(po0622),
    .po0623(po0623),
    .po0624(po0624),
    .po0625(po0625),
    .po0626(po0626),
    .po0627(po0627),
    .po0628(po0628),
    .po0629(po0629),
    .po0630(po0630),
    .po0631(po0631),
    .po0632(po0632),
    .po0633(po0633),
    .po0634(po0634),
    .po0635(po0635),
    .po0636(po0636),
    .po0637(po0637),
    .po0638(po0638),
    .po0639(po0639),
    .po0640(po0640),
    .po0641(po0641),
    .po0642(po0642),
    .po0643(po0643),
    .po0644(po0644),
    .po0645(po0645),
    .po0646(po0646),
    .po0647(po0647),
    .po0648(po0648),
    .po0649(po0649),
    .po0650(po0650),
    .po0651(po0651),
    .po0652(po0652),
    .po0653(po0653),
    .po0654(po0654),
    .po0655(po0655),
    .po0656(po0656),
    .po0657(po0657),
    .po0658(po0658),
    .po0659(po0659),
    .po0660(po0660),
    .po0661(po0661),
    .po0662(po0662),
    .po0663(po0663),
    .po0664(po0664),
    .po0665(po0665),
    .po0666(po0666),
    .po0667(po0667),
    .po0668(po0668),
    .po0669(po0669),
    .po0670(po0670),
    .po0671(po0671),
    .po0672(po0672),
    .po0673(po0673),
    .po0674(po0674),
    .po0675(po0675),
    .po0676(po0676),
    .po0677(po0677),
    .po0678(po0678),
    .po0679(po0679),
    .po0680(po0680),
    .po0681(po0681),
    .po0682(po0682),
    .po0683(po0683),
    .po0684(po0684),
    .po0685(po0685),
    .po0686(po0686),
    .po0687(po0687),
    .po0688(po0688),
    .po0689(po0689),
    .po0690(po0690),
    .po0691(po0691),
    .po0692(po0692),
    .po0693(po0693),
    .po0694(po0694),
    .po0695(po0695),
    .po0696(po0696),
    .po0697(po0697),
    .po0698(po0698),
    .po0699(po0699),
    .po0700(po0700),
    .po0701(po0701),
    .po0702(po0702),
    .po0703(po0703),
    .po0704(po0704),
    .po0705(po0705),
    .po0706(po0706),
    .po0707(po0707),
    .po0708(po0708),
    .po0709(po0709),
    .po0710(po0710),
    .po0711(po0711),
    .po0712(po0712),
    .po0713(po0713),
    .po0714(po0714),
    .po0715(po0715),
    .po0716(po0716),
    .po0717(po0717),
    .po0718(po0718),
    .po0719(po0719),
    .po0720(po0720),
    .po0721(po0721),
    .po0722(po0722),
    .po0723(po0723),
    .po0724(po0724),
    .po0725(po0725),
    .po0726(po0726),
    .po0727(po0727),
    .po0728(po0728),
    .po0729(po0729),
    .po0730(po0730),
    .po0731(po0731),
    .po0732(po0732),
    .po0733(po0733),
    .po0734(po0734),
    .po0735(po0735),
    .po0736(po0736),
    .po0737(po0737),
    .po0738(po0738),
    .po0739(po0739),
    .po0740(po0740),
    .po0741(po0741),
    .po0742(po0742),
    .po0743(po0743),
    .po0744(po0744),
    .po0745(po0745),
    .po0746(po0746),
    .po0747(po0747),
    .po0748(po0748),
    .po0749(po0749),
    .po0750(po0750),
    .po0751(po0751),
    .po0752(po0752),
    .po0753(po0753),
    .po0754(po0754),
    .po0755(po0755),
    .po0756(po0756),
    .po0757(po0757),
    .po0758(po0758),
    .po0759(po0759),
    .po0760(po0760),
    .po0761(po0761),
    .po0762(po0762),
    .po0763(po0763),
    .po0764(po0764),
    .po0765(po0765),
    .po0766(po0766),
    .po0767(po0767),
    .po0768(po0768),
    .po0769(po0769),
    .po0770(po0770),
    .po0771(po0771),
    .po0772(po0772),
    .po0773(po0773),
    .po0774(po0774),
    .po0775(po0775),
    .po0776(po0776),
    .po0777(po0777),
    .po0778(po0778),
    .po0779(po0779),
    .po0780(po0780),
    .po0781(po0781),
    .po0782(po0782),
    .po0783(po0783),
    .po0784(po0784),
    .po0785(po0785),
    .po0786(po0786),
    .po0787(po0787),
    .po0788(po0788),
    .po0789(po0789),
    .po0790(po0790),
    .po0791(po0791),
    .po0792(po0792),
    .po0793(po0793),
    .po0794(po0794),
    .po0795(po0795),
    .po0796(po0796),
    .po0797(po0797),
    .po0798(po0798),
    .po0799(po0799),
    .po0800(po0800),
    .po0801(po0801),
    .po0802(po0802),
    .po0803(po0803),
    .po0804(po0804),
    .po0805(po0805),
    .po0806(po0806),
    .po0807(po0807),
    .po0808(po0808),
    .po0809(po0809),
    .po0810(po0810),
    .po0811(po0811),
    .po0812(po0812),
    .po0813(po0813),
    .po0814(po0814),
    .po0815(po0815),
    .po0816(po0816),
    .po0817(po0817),
    .po0818(po0818),
    .po0819(po0819),
    .po0820(po0820),
    .po0821(po0821),
    .po0822(po0822),
    .po0823(po0823),
    .po0824(po0824),
    .po0825(po0825),
    .po0826(po0826),
    .po0827(po0827),
    .po0828(po0828),
    .po0829(po0829),
    .po0830(po0830),
    .po0831(po0831),
    .po0832(po0832),
    .po0833(po0833),
    .po0834(po0834),
    .po0835(po0835),
    .po0836(po0836),
    .po0837(po0837),
    .po0838(po0838),
    .po0839(po0839),
    .po0840(po0840),
    .po0841(po0841),
    .po0842(po0842),
    .po0843(po0843),
    .po0844(po0844),
    .po0845(po0845),
    .po0846(po0846),
    .po0847(po0847),
    .po0848(po0848),
    .po0849(po0849),
    .po0850(po0850),
    .po0851(po0851),
    .po0852(po0852),
    .po0853(po0853),
    .po0854(po0854),
    .po0855(po0855),
    .po0856(po0856),
    .po0857(po0857),
    .po0858(po0858),
    .po0859(po0859),
    .po0860(po0860),
    .po0861(po0861),
    .po0862(po0862),
    .po0863(po0863),
    .po0864(po0864),
    .po0865(po0865),
    .po0866(po0866),
    .po0867(po0867),
    .po0868(po0868),
    .po0869(po0869),
    .po0870(po0870),
    .po0871(po0871),
    .po0872(po0872),
    .po0873(po0873),
    .po0874(po0874),
    .po0875(po0875),
    .po0876(po0876),
    .po0877(po0877),
    .po0878(po0878),
    .po0879(po0879),
    .po0880(po0880),
    .po0881(po0881),
    .po0882(po0882),
    .po0883(po0883),
    .po0884(po0884),
    .po0885(po0885),
    .po0886(po0886),
    .po0887(po0887),
    .po0888(po0888),
    .po0889(po0889),
    .po0890(po0890),
    .po0891(po0891),
    .po0892(po0892),
    .po0893(po0893),
    .po0894(po0894),
    .po0895(po0895),
    .po0896(po0896),
    .po0897(po0897),
    .po0898(po0898),
    .po0899(po0899),
    .po0900(po0900),
    .po0901(po0901),
    .po0902(po0902),
    .po0903(po0903),
    .po0904(po0904),
    .po0905(po0905),
    .po0906(po0906),
    .po0907(po0907),
    .po0908(po0908),
    .po0909(po0909),
    .po0910(po0910),
    .po0911(po0911),
    .po0912(po0912),
    .po0913(po0913),
    .po0914(po0914),
    .po0915(po0915),
    .po0916(po0916),
    .po0917(po0917),
    .po0918(po0918),
    .po0919(po0919),
    .po0920(po0920),
    .po0921(po0921),
    .po0922(po0922),
    .po0923(po0923),
    .po0924(po0924),
    .po0925(po0925),
    .po0926(po0926),
    .po0927(po0927),
    .po0928(po0928),
    .po0929(po0929),
    .po0930(po0930),
    .po0931(po0931),
    .po0932(po0932),
    .po0933(po0933),
    .po0934(po0934),
    .po0935(po0935),
    .po0936(po0936),
    .po0937(po0937),
    .po0938(po0938),
    .po0939(po0939),
    .po0940(po0940),
    .po0941(po0941),
    .po0942(po0942),
    .po0943(po0943),
    .po0944(po0944),
    .po0945(po0945),
    .po0946(po0946),
    .po0947(po0947),
    .po0948(po0948),
    .po0949(po0949),
    .po0950(po0950),
    .po0951(po0951),
    .po0952(po0952),
    .po0953(po0953),
    .po0954(po0954),
    .po0955(po0955),
    .po0956(po0956),
    .po0957(po0957),
    .po0958(po0958),
    .po0959(po0959),
    .po0960(po0960),
    .po0961(po0961),
    .po0962(po0962),
    .po0963(po0963),
    .po0964(po0964),
    .po0965(po0965),
    .po0966(po0966),
    .po0967(po0967),
    .po0968(po0968),
    .po0969(po0969),
    .po0970(po0970),
    .po0971(po0971),
    .po0972(po0972),
    .po0973(po0973),
    .po0974(po0974),
    .po0975(po0975),
    .po0976(po0976),
    .po0977(po0977),
    .po0978(po0978),
    .po0979(po0979),
    .po0980(po0980),
    .po0981(po0981),
    .po0982(po0982),
    .po0983(po0983),
    .po0984(po0984),
    .po0985(po0985),
    .po0986(po0986),
    .po0987(po0987),
    .po0988(po0988),
    .po0989(po0989),
    .po0990(po0990),
    .po0991(po0991),
    .po0992(po0992),
    .po0993(po0993),
    .po0994(po0994),
    .po0995(po0995),
    .po0996(po0996),
    .po0997(po0997),
    .po0998(po0998),
    .po0999(po0999),
    .po1000(po1000),
    .po1001(po1001),
    .po1002(po1002),
    .po1003(po1003),
    .po1004(po1004),
    .po1005(po1005),
    .po1006(po1006),
    .po1007(po1007),
    .po1008(po1008),
    .po1009(po1009),
    .po1010(po1010),
    .po1011(po1011),
    .po1012(po1012),
    .po1013(po1013),
    .po1014(po1014),
    .po1015(po1015),
    .po1016(po1016),
    .po1017(po1017),
    .po1018(po1018),
    .po1019(po1019),
    .po1020(po1020),
    .po1021(po1021),
    .po1022(po1022),
    .po1023(po1023),
    .po1024(po1024),
    .po1025(po1025),
    .po1026(po1026),
    .po1027(po1027),
    .po1028(po1028),
    .po1029(po1029),
    .po1030(po1030),
    .po1031(po1031),
    .po1032(po1032),
    .po1033(po1033),
    .po1034(po1034),
    .po1035(po1035),
    .po1036(po1036),
    .po1037(po1037),
    .po1038(po1038),
    .po1039(po1039),
    .po1040(po1040),
    .po1041(po1041),
    .po1042(po1042),
    .po1043(po1043),
    .po1044(po1044),
    .po1045(po1045),
    .po1046(po1046),
    .po1047(po1047),
    .po1048(po1048),
    .po1049(po1049),
    .po1050(po1050),
    .po1051(po1051),
    .po1052(po1052),
    .po1053(po1053),
    .po1054(po1054),
    .po1055(po1055),
    .po1056(po1056),
    .po1057(po1057),
    .po1058(po1058),
    .po1059(po1059),
    .po1060(po1060),
    .po1061(po1061),
    .po1062(po1062),
    .po1063(po1063),
    .po1064(po1064),
    .po1065(po1065),
    .po1066(po1066),
    .po1067(po1067),
    .po1068(po1068),
    .po1069(po1069),
    .po1070(po1070),
    .po1071(po1071),
    .po1072(po1072),
    .po1073(po1073),
    .po1074(po1074),
    .po1075(po1075),
    .po1076(po1076),
    .po1077(po1077),
    .po1078(po1078),
    .po1079(po1079),
    .po1080(po1080),
    .po1081(po1081),
    .po1082(po1082),
    .po1083(po1083),
    .po1084(po1084),
    .po1085(po1085),
    .po1086(po1086),
    .po1087(po1087),
    .po1088(po1088),
    .po1089(po1089),
    .po1090(po1090),
    .po1091(po1091),
    .po1092(po1092),
    .po1093(po1093),
    .po1094(po1094),
    .po1095(po1095),
    .po1096(po1096),
    .po1097(po1097),
    .po1098(po1098),
    .po1099(po1099),
    .po1100(po1100),
    .po1101(po1101),
    .po1102(po1102),
    .po1103(po1103),
    .po1104(po1104),
    .po1105(po1105),
    .po1106(po1106),
    .po1107(po1107),
    .po1108(po1108),
    .po1109(po1109),
    .po1110(po1110),
    .po1111(po1111),
    .po1112(po1112),
    .po1113(po1113),
    .po1114(po1114),
    .po1115(po1115),
    .po1116(po1116),
    .po1117(po1117),
    .po1118(po1118),
    .po1119(po1119),
    .po1120(po1120),
    .po1121(po1121),
    .po1122(po1122),
    .po1123(po1123),
    .po1124(po1124),
    .po1125(po1125),
    .po1126(po1126),
    .po1127(po1127),
    .po1128(po1128),
    .po1129(po1129),
    .po1130(po1130),
    .po1131(po1131),
    .po1132(po1132),
    .po1133(po1133),
    .po1134(po1134),
    .po1135(po1135),
    .po1136(po1136),
    .po1137(po1137),
    .po1138(po1138),
    .po1139(po1139),
    .po1140(po1140),
    .po1141(po1141),
    .po1142(po1142),
    .po1143(po1143),
    .po1144(po1144),
    .po1145(po1145),
    .po1146(po1146),
    .po1147(po1147),
    .po1148(po1148),
    .po1149(po1149),
    .po1150(po1150),
    .po1151(po1151),
    .po1152(po1152),
    .po1153(po1153),
    .po1154(po1154),
    .po1155(po1155),
    .po1156(po1156),
    .po1157(po1157),
    .po1158(po1158),
    .po1159(po1159),
    .po1160(po1160),
    .po1161(po1161),
    .po1162(po1162),
    .po1163(po1163),
    .po1164(po1164),
    .po1165(po1165),
    .po1166(po1166),
    .po1167(po1167),
    .po1168(po1168),
    .po1169(po1169),
    .po1170(po1170),
    .po1171(po1171),
    .po1172(po1172),
    .po1173(po1173),
    .po1174(po1174),
    .po1175(po1175),
    .po1176(po1176),
    .po1177(po1177),
    .po1178(po1178),
    .po1179(po1179),
    .po1180(po1180),
    .po1181(po1181),
    .po1182(po1182),
    .po1183(po1183),
    .po1184(po1184),
    .po1185(po1185),
    .po1186(po1186),
    .po1187(po1187),
    .po1188(po1188),
    .po1189(po1189),
    .po1190(po1190),
    .po1191(po1191),
    .po1192(po1192),
    .po1193(po1193),
    .po1194(po1194),
    .po1195(po1195),
    .po1196(po1196),
    .po1197(po1197),
    .po1198(po1198),
    .po1199(po1199),
    .po1200(po1200),
    .po1201(po1201),
    .po1202(po1202),
    .po1203(po1203),
    .po1204(po1204),
    .po1205(po1205),
    .po1206(po1206),
    .po1207(po1207),
    .po1208(po1208),
    .po1209(po1209),
    .po1210(po1210),
    .po1211(po1211),
    .po1212(po1212),
    .po1213(po1213),
    .po1214(po1214),
    .po1215(po1215),
    .po1216(po1216),
    .po1217(po1217),
    .po1218(po1218),
    .po1219(po1219),
    .po1220(po1220),
    .po1221(po1221),
    .po1222(po1222),
    .po1223(po1223),
    .po1224(po1224),
    .po1225(po1225),
    .po1226(po1226),
    .po1227(po1227),
    .po1228(po1228),
    .po1229(po1229),
    .po1230(po1230)
  );

  // Random function
  integer SEED = 6;
  function [7:0] urand(input integer s);
    urand = $random(s) & 8'hFF;
  endfunction

  // Main stimulus (combinational)
  integer i;
  parameter CYCLES = 512;
  parameter PRINT_EVERY = 1;

  initial begin
    pi0000= 0;
    pi0001= 0;
    pi0002= 0;
    pi0003= 0;
    pi0004= 0;
    pi0005= 0;
    pi0006= 0;
    pi0007= 0;
    pi0008= 0;
    pi0009= 0;
    pi0010= 0;
    pi0011= 0;
    pi0012= 0;
    pi0013= 0;
    pi0014= 0;
    pi0015= 0;
    pi0016= 0;
    pi0017= 0;
    pi0018= 0;
    pi0019= 0;
    pi0020= 0;
    pi0021= 0;
    pi0022= 0;
    pi0023= 0;
    pi0024= 0;
    pi0025= 0;
    pi0026= 0;
    pi0027= 0;
    pi0028= 0;
    pi0029= 0;
    pi0030= 0;
    pi0031= 0;
    pi0032= 0;
    pi0033= 0;
    pi0034= 0;
    pi0035= 0;
    pi0036= 0;
    pi0037= 0;
    pi0038= 0;
    pi0039= 0;
    pi0040= 0;
    pi0041= 0;
    pi0042= 0;
    pi0043= 0;
    pi0044= 0;
    pi0045= 0;
    pi0046= 0;
    pi0047= 0;
    pi0048= 0;
    pi0049= 0;
    pi0050= 0;
    pi0051= 0;
    pi0052= 0;
    pi0053= 0;
    pi0054= 0;
    pi0055= 0;
    pi0056= 0;
    pi0057= 0;
    pi0058= 0;
    pi0059= 0;
    pi0060= 0;
    pi0061= 0;
    pi0062= 0;
    pi0063= 0;
    pi0064= 0;
    pi0065= 0;
    pi0066= 0;
    pi0067= 0;
    pi0068= 0;
    pi0069= 0;
    pi0070= 0;
    pi0071= 0;
    pi0072= 0;
    pi0073= 0;
    pi0074= 0;
    pi0075= 0;
    pi0076= 0;
    pi0077= 0;
    pi0078= 0;
    pi0079= 0;
    pi0080= 0;
    pi0081= 0;
    pi0082= 0;
    pi0083= 0;
    pi0084= 0;
    pi0085= 0;
    pi0086= 0;
    pi0087= 0;
    pi0088= 0;
    pi0089= 0;
    pi0090= 0;
    pi0091= 0;
    pi0092= 0;
    pi0093= 0;
    pi0094= 0;
    pi0095= 0;
    pi0096= 0;
    pi0097= 0;
    pi0098= 0;
    pi0099= 0;
    pi0100= 0;
    pi0101= 0;
    pi0102= 0;
    pi0103= 0;
    pi0104= 0;
    pi0105= 0;
    pi0106= 0;
    pi0107= 0;
    pi0108= 0;
    pi0109= 0;
    pi0110= 0;
    pi0111= 0;
    pi0112= 0;
    pi0113= 0;
    pi0114= 0;
    pi0115= 0;
    pi0116= 0;
    pi0117= 0;
    pi0118= 0;
    pi0119= 0;
    pi0120= 0;
    pi0121= 0;
    pi0122= 0;
    pi0123= 0;
    pi0124= 0;
    pi0125= 0;
    pi0126= 0;
    pi0127= 0;
    pi0128= 0;
    pi0129= 0;
    pi0130= 0;
    pi0131= 0;
    pi0132= 0;
    pi0133= 0;
    pi0134= 0;
    pi0135= 0;
    pi0136= 0;
    pi0137= 0;
    pi0138= 0;
    pi0139= 0;
    pi0140= 0;
    pi0141= 0;
    pi0142= 0;
    pi0143= 0;
    pi0144= 0;
    pi0145= 0;
    pi0146= 0;
    pi0147= 0;
    pi0148= 0;
    pi0149= 0;
    pi0150= 0;
    pi0151= 0;
    pi0152= 0;
    pi0153= 0;
    pi0154= 0;
    pi0155= 0;
    pi0156= 0;
    pi0157= 0;
    pi0158= 0;
    pi0159= 0;
    pi0160= 0;
    pi0161= 0;
    pi0162= 0;
    pi0163= 0;
    pi0164= 0;
    pi0165= 0;
    pi0166= 0;
    pi0167= 0;
    pi0168= 0;
    pi0169= 0;
    pi0170= 0;
    pi0171= 0;
    pi0172= 0;
    pi0173= 0;
    pi0174= 0;
    pi0175= 0;
    pi0176= 0;
    pi0177= 0;
    pi0178= 0;
    pi0179= 0;
    pi0180= 0;
    pi0181= 0;
    pi0182= 0;
    pi0183= 0;
    pi0184= 0;
    pi0185= 0;
    pi0186= 0;
    pi0187= 0;
    pi0188= 0;
    pi0189= 0;
    pi0190= 0;
    pi0191= 0;
    pi0192= 0;
    pi0193= 0;
    pi0194= 0;
    pi0195= 0;
    pi0196= 0;
    pi0197= 0;
    pi0198= 0;
    pi0199= 0;
    pi0200= 0;
    pi0201= 0;
    pi0202= 0;
    pi0203= 0;
    pi0204= 0;
    pi0205= 0;
    pi0206= 0;
    pi0207= 0;
    pi0208= 0;
    pi0209= 0;
    pi0210= 0;
    pi0211= 0;
    pi0212= 0;
    pi0213= 0;
    pi0214= 0;
    pi0215= 0;
    pi0216= 0;
    pi0217= 0;
    pi0218= 0;
    pi0219= 0;
    pi0220= 0;
    pi0221= 0;
    pi0222= 0;
    pi0223= 0;
    pi0224= 0;
    pi0225= 0;
    pi0226= 0;
    pi0227= 0;
    pi0228= 0;
    pi0229= 0;
    pi0230= 0;
    pi0231= 0;
    pi0232= 0;
    pi0233= 0;
    pi0234= 0;
    pi0235= 0;
    pi0236= 0;
    pi0237= 0;
    pi0238= 0;
    pi0239= 0;
    pi0240= 0;
    pi0241= 0;
    pi0242= 0;
    pi0243= 0;
    pi0244= 0;
    pi0245= 0;
    pi0246= 0;
    pi0247= 0;
    pi0248= 0;
    pi0249= 0;
    pi0250= 0;
    pi0251= 0;
    pi0252= 0;
    pi0253= 0;
    pi0254= 0;
    pi0255= 0;
    pi0256= 0;
    pi0257= 0;
    pi0258= 0;
    pi0259= 0;
    pi0260= 0;
    pi0261= 0;
    pi0262= 0;
    pi0263= 0;
    pi0264= 0;
    pi0265= 0;
    pi0266= 0;
    pi0267= 0;
    pi0268= 0;
    pi0269= 0;
    pi0270= 0;
    pi0271= 0;
    pi0272= 0;
    pi0273= 0;
    pi0274= 0;
    pi0275= 0;
    pi0276= 0;
    pi0277= 0;
    pi0278= 0;
    pi0279= 0;
    pi0280= 0;
    pi0281= 0;
    pi0282= 0;
    pi0283= 0;
    pi0284= 0;
    pi0285= 0;
    pi0286= 0;
    pi0287= 0;
    pi0288= 0;
    pi0289= 0;
    pi0290= 0;
    pi0291= 0;
    pi0292= 0;
    pi0293= 0;
    pi0294= 0;
    pi0295= 0;
    pi0296= 0;
    pi0297= 0;
    pi0298= 0;
    pi0299= 0;
    pi0300= 0;
    pi0301= 0;
    pi0302= 0;
    pi0303= 0;
    pi0304= 0;
    pi0305= 0;
    pi0306= 0;
    pi0307= 0;
    pi0308= 0;
    pi0309= 0;
    pi0310= 0;
    pi0311= 0;
    pi0312= 0;
    pi0313= 0;
    pi0314= 0;
    pi0315= 0;
    pi0316= 0;
    pi0317= 0;
    pi0318= 0;
    pi0319= 0;
    pi0320= 0;
    pi0321= 0;
    pi0322= 0;
    pi0323= 0;
    pi0324= 0;
    pi0325= 0;
    pi0326= 0;
    pi0327= 0;
    pi0328= 0;
    pi0329= 0;
    pi0330= 0;
    pi0331= 0;
    pi0332= 0;
    pi0333= 0;
    pi0334= 0;
    pi0335= 0;
    pi0336= 0;
    pi0337= 0;
    pi0338= 0;
    pi0339= 0;
    pi0340= 0;
    pi0341= 0;
    pi0342= 0;
    pi0343= 0;
    pi0344= 0;
    pi0345= 0;
    pi0346= 0;
    pi0347= 0;
    pi0348= 0;
    pi0349= 0;
    pi0350= 0;
    pi0351= 0;
    pi0352= 0;
    pi0353= 0;
    pi0354= 0;
    pi0355= 0;
    pi0356= 0;
    pi0357= 0;
    pi0358= 0;
    pi0359= 0;
    pi0360= 0;
    pi0361= 0;
    pi0362= 0;
    pi0363= 0;
    pi0364= 0;
    pi0365= 0;
    pi0366= 0;
    pi0367= 0;
    pi0368= 0;
    pi0369= 0;
    pi0370= 0;
    pi0371= 0;
    pi0372= 0;
    pi0373= 0;
    pi0374= 0;
    pi0375= 0;
    pi0376= 0;
    pi0377= 0;
    pi0378= 0;
    pi0379= 0;
    pi0380= 0;
    pi0381= 0;
    pi0382= 0;
    pi0383= 0;
    pi0384= 0;
    pi0385= 0;
    pi0386= 0;
    pi0387= 0;
    pi0388= 0;
    pi0389= 0;
    pi0390= 0;
    pi0391= 0;
    pi0392= 0;
    pi0393= 0;
    pi0394= 0;
    pi0395= 0;
    pi0396= 0;
    pi0397= 0;
    pi0398= 0;
    pi0399= 0;
    pi0400= 0;
    pi0401= 0;
    pi0402= 0;
    pi0403= 0;
    pi0404= 0;
    pi0405= 0;
    pi0406= 0;
    pi0407= 0;
    pi0408= 0;
    pi0409= 0;
    pi0410= 0;
    pi0411= 0;
    pi0412= 0;
    pi0413= 0;
    pi0414= 0;
    pi0415= 0;
    pi0416= 0;
    pi0417= 0;
    pi0418= 0;
    pi0419= 0;
    pi0420= 0;
    pi0421= 0;
    pi0422= 0;
    pi0423= 0;
    pi0424= 0;
    pi0425= 0;
    pi0426= 0;
    pi0427= 0;
    pi0428= 0;
    pi0429= 0;
    pi0430= 0;
    pi0431= 0;
    pi0432= 0;
    pi0433= 0;
    pi0434= 0;
    pi0435= 0;
    pi0436= 0;
    pi0437= 0;
    pi0438= 0;
    pi0439= 0;
    pi0440= 0;
    pi0441= 0;
    pi0442= 0;
    pi0443= 0;
    pi0444= 0;
    pi0445= 0;
    pi0446= 0;
    pi0447= 0;
    pi0448= 0;
    pi0449= 0;
    pi0450= 0;
    pi0451= 0;
    pi0452= 0;
    pi0453= 0;
    pi0454= 0;
    pi0455= 0;
    pi0456= 0;
    pi0457= 0;
    pi0458= 0;
    pi0459= 0;
    pi0460= 0;
    pi0461= 0;
    pi0462= 0;
    pi0463= 0;
    pi0464= 0;
    pi0465= 0;
    pi0466= 0;
    pi0467= 0;
    pi0468= 0;
    pi0469= 0;
    pi0470= 0;
    pi0471= 0;
    pi0472= 0;
    pi0473= 0;
    pi0474= 0;
    pi0475= 0;
    pi0476= 0;
    pi0477= 0;
    pi0478= 0;
    pi0479= 0;
    pi0480= 0;
    pi0481= 0;
    pi0482= 0;
    pi0483= 0;
    pi0484= 0;
    pi0485= 0;
    pi0486= 0;
    pi0487= 0;
    pi0488= 0;
    pi0489= 0;
    pi0490= 0;
    pi0491= 0;
    pi0492= 0;
    pi0493= 0;
    pi0494= 0;
    pi0495= 0;
    pi0496= 0;
    pi0497= 0;
    pi0498= 0;
    pi0499= 0;
    pi0500= 0;
    pi0501= 0;
    pi0502= 0;
    pi0503= 0;
    pi0504= 0;
    pi0505= 0;
    pi0506= 0;
    pi0507= 0;
    pi0508= 0;
    pi0509= 0;
    pi0510= 0;
    pi0511= 0;
    pi0512= 0;
    pi0513= 0;
    pi0514= 0;
    pi0515= 0;
    pi0516= 0;
    pi0517= 0;
    pi0518= 0;
    pi0519= 0;
    pi0520= 0;
    pi0521= 0;
    pi0522= 0;
    pi0523= 0;
    pi0524= 0;
    pi0525= 0;
    pi0526= 0;
    pi0527= 0;
    pi0528= 0;
    pi0529= 0;
    pi0530= 0;
    pi0531= 0;
    pi0532= 0;
    pi0533= 0;
    pi0534= 0;
    pi0535= 0;
    pi0536= 0;
    pi0537= 0;
    pi0538= 0;
    pi0539= 0;
    pi0540= 0;
    pi0541= 0;
    pi0542= 0;
    pi0543= 0;
    pi0544= 0;
    pi0545= 0;
    pi0546= 0;
    pi0547= 0;
    pi0548= 0;
    pi0549= 0;
    pi0550= 0;
    pi0551= 0;
    pi0552= 0;
    pi0553= 0;
    pi0554= 0;
    pi0555= 0;
    pi0556= 0;
    pi0557= 0;
    pi0558= 0;
    pi0559= 0;
    pi0560= 0;
    pi0561= 0;
    pi0562= 0;
    pi0563= 0;
    pi0564= 0;
    pi0565= 0;
    pi0566= 0;
    pi0567= 0;
    pi0568= 0;
    pi0569= 0;
    pi0570= 0;
    pi0571= 0;
    pi0572= 0;
    pi0573= 0;
    pi0574= 0;
    pi0575= 0;
    pi0576= 0;
    pi0577= 0;
    pi0578= 0;
    pi0579= 0;
    pi0580= 0;
    pi0581= 0;
    pi0582= 0;
    pi0583= 0;
    pi0584= 0;
    pi0585= 0;
    pi0586= 0;
    pi0587= 0;
    pi0588= 0;
    pi0589= 0;
    pi0590= 0;
    pi0591= 0;
    pi0592= 0;
    pi0593= 0;
    pi0594= 0;
    pi0595= 0;
    pi0596= 0;
    pi0597= 0;
    pi0598= 0;
    pi0599= 0;
    pi0600= 0;
    pi0601= 0;
    pi0602= 0;
    pi0603= 0;
    pi0604= 0;
    pi0605= 0;
    pi0606= 0;
    pi0607= 0;
    pi0608= 0;
    pi0609= 0;
    pi0610= 0;
    pi0611= 0;
    pi0612= 0;
    pi0613= 0;
    pi0614= 0;
    pi0615= 0;
    pi0616= 0;
    pi0617= 0;
    pi0618= 0;
    pi0619= 0;
    pi0620= 0;
    pi0621= 0;
    pi0622= 0;
    pi0623= 0;
    pi0624= 0;
    pi0625= 0;
    pi0626= 0;
    pi0627= 0;
    pi0628= 0;
    pi0629= 0;
    pi0630= 0;
    pi0631= 0;
    pi0632= 0;
    pi0633= 0;
    pi0634= 0;
    pi0635= 0;
    pi0636= 0;
    pi0637= 0;
    pi0638= 0;
    pi0639= 0;
    pi0640= 0;
    pi0641= 0;
    pi0642= 0;
    pi0643= 0;
    pi0644= 0;
    pi0645= 0;
    pi0646= 0;
    pi0647= 0;
    pi0648= 0;
    pi0649= 0;
    pi0650= 0;
    pi0651= 0;
    pi0652= 0;
    pi0653= 0;
    pi0654= 0;
    pi0655= 0;
    pi0656= 0;
    pi0657= 0;
    pi0658= 0;
    pi0659= 0;
    pi0660= 0;
    pi0661= 0;
    pi0662= 0;
    pi0663= 0;
    pi0664= 0;
    pi0665= 0;
    pi0666= 0;
    pi0667= 0;
    pi0668= 0;
    pi0669= 0;
    pi0670= 0;
    pi0671= 0;
    pi0672= 0;
    pi0673= 0;
    pi0674= 0;
    pi0675= 0;
    pi0676= 0;
    pi0677= 0;
    pi0678= 0;
    pi0679= 0;
    pi0680= 0;
    pi0681= 0;
    pi0682= 0;
    pi0683= 0;
    pi0684= 0;
    pi0685= 0;
    pi0686= 0;
    pi0687= 0;
    pi0688= 0;
    pi0689= 0;
    pi0690= 0;
    pi0691= 0;
    pi0692= 0;
    pi0693= 0;
    pi0694= 0;
    pi0695= 0;
    pi0696= 0;
    pi0697= 0;
    pi0698= 0;
    pi0699= 0;
    pi0700= 0;
    pi0701= 0;
    pi0702= 0;
    pi0703= 0;
    pi0704= 0;
    pi0705= 0;
    pi0706= 0;
    pi0707= 0;
    pi0708= 0;
    pi0709= 0;
    pi0710= 0;
    pi0711= 0;
    pi0712= 0;
    pi0713= 0;
    pi0714= 0;
    pi0715= 0;
    pi0716= 0;
    pi0717= 0;
    pi0718= 0;
    pi0719= 0;
    pi0720= 0;
    pi0721= 0;
    pi0722= 0;
    pi0723= 0;
    pi0724= 0;
    pi0725= 0;
    pi0726= 0;
    pi0727= 0;
    pi0728= 0;
    pi0729= 0;
    pi0730= 0;
    pi0731= 0;
    pi0732= 0;
    pi0733= 0;
    pi0734= 0;
    pi0735= 0;
    pi0736= 0;
    pi0737= 0;
    pi0738= 0;
    pi0739= 0;
    pi0740= 0;
    pi0741= 0;
    pi0742= 0;
    pi0743= 0;
    pi0744= 0;
    pi0745= 0;
    pi0746= 0;
    pi0747= 0;
    pi0748= 0;
    pi0749= 0;
    pi0750= 0;
    pi0751= 0;
    pi0752= 0;
    pi0753= 0;
    pi0754= 0;
    pi0755= 0;
    pi0756= 0;
    pi0757= 0;
    pi0758= 0;
    pi0759= 0;
    pi0760= 0;
    pi0761= 0;
    pi0762= 0;
    pi0763= 0;
    pi0764= 0;
    pi0765= 0;
    pi0766= 0;
    pi0767= 0;
    pi0768= 0;
    pi0769= 0;
    pi0770= 0;
    pi0771= 0;
    pi0772= 0;
    pi0773= 0;
    pi0774= 0;
    pi0775= 0;
    pi0776= 0;
    pi0777= 0;
    pi0778= 0;
    pi0779= 0;
    pi0780= 0;
    pi0781= 0;
    pi0782= 0;
    pi0783= 0;
    pi0784= 0;
    pi0785= 0;
    pi0786= 0;
    pi0787= 0;
    pi0788= 0;
    pi0789= 0;
    pi0790= 0;
    pi0791= 0;
    pi0792= 0;
    pi0793= 0;
    pi0794= 0;
    pi0795= 0;
    pi0796= 0;
    pi0797= 0;
    pi0798= 0;
    pi0799= 0;
    pi0800= 0;
    pi0801= 0;
    pi0802= 0;
    pi0803= 0;
    pi0804= 0;
    pi0805= 0;
    pi0806= 0;
    pi0807= 0;
    pi0808= 0;
    pi0809= 0;
    pi0810= 0;
    pi0811= 0;
    pi0812= 0;
    pi0813= 0;
    pi0814= 0;
    pi0815= 0;
    pi0816= 0;
    pi0817= 0;
    pi0818= 0;
    pi0819= 0;
    pi0820= 0;
    pi0821= 0;
    pi0822= 0;
    pi0823= 0;
    pi0824= 0;
    pi0825= 0;
    pi0826= 0;
    pi0827= 0;
    pi0828= 0;
    pi0829= 0;
    pi0830= 0;
    pi0831= 0;
    pi0832= 0;
    pi0833= 0;
    pi0834= 0;
    pi0835= 0;
    pi0836= 0;
    pi0837= 0;
    pi0838= 0;
    pi0839= 0;
    pi0840= 0;
    pi0841= 0;
    pi0842= 0;
    pi0843= 0;
    pi0844= 0;
    pi0845= 0;
    pi0846= 0;
    pi0847= 0;
    pi0848= 0;
    pi0849= 0;
    pi0850= 0;
    pi0851= 0;
    pi0852= 0;
    pi0853= 0;
    pi0854= 0;
    pi0855= 0;
    pi0856= 0;
    pi0857= 0;
    pi0858= 0;
    pi0859= 0;
    pi0860= 0;
    pi0861= 0;
    pi0862= 0;
    pi0863= 0;
    pi0864= 0;
    pi0865= 0;
    pi0866= 0;
    pi0867= 0;
    pi0868= 0;
    pi0869= 0;
    pi0870= 0;
    pi0871= 0;
    pi0872= 0;
    pi0873= 0;
    pi0874= 0;
    pi0875= 0;
    pi0876= 0;
    pi0877= 0;
    pi0878= 0;
    pi0879= 0;
    pi0880= 0;
    pi0881= 0;
    pi0882= 0;
    pi0883= 0;
    pi0884= 0;
    pi0885= 0;
    pi0886= 0;
    pi0887= 0;
    pi0888= 0;
    pi0889= 0;
    pi0890= 0;
    pi0891= 0;
    pi0892= 0;
    pi0893= 0;
    pi0894= 0;
    pi0895= 0;
    pi0896= 0;
    pi0897= 0;
    pi0898= 0;
    pi0899= 0;
    pi0900= 0;
    pi0901= 0;
    pi0902= 0;
    pi0903= 0;
    pi0904= 0;
    pi0905= 0;
    pi0906= 0;
    pi0907= 0;
    pi0908= 0;
    pi0909= 0;
    pi0910= 0;
    pi0911= 0;
    pi0912= 0;
    pi0913= 0;
    pi0914= 0;
    pi0915= 0;
    pi0916= 0;
    pi0917= 0;
    pi0918= 0;
    pi0919= 0;
    pi0920= 0;
    pi0921= 0;
    pi0922= 0;
    pi0923= 0;
    pi0924= 0;
    pi0925= 0;
    pi0926= 0;
    pi0927= 0;
    pi0928= 0;
    pi0929= 0;
    pi0930= 0;
    pi0931= 0;
    pi0932= 0;
    pi0933= 0;
    pi0934= 0;
    pi0935= 0;
    pi0936= 0;
    pi0937= 0;
    pi0938= 0;
    pi0939= 0;
    pi0940= 0;
    pi0941= 0;
    pi0942= 0;
    pi0943= 0;
    pi0944= 0;
    pi0945= 0;
    pi0946= 0;
    pi0947= 0;
    pi0948= 0;
    pi0949= 0;
    pi0950= 0;
    pi0951= 0;
    pi0952= 0;
    pi0953= 0;
    pi0954= 0;
    pi0955= 0;
    pi0956= 0;
    pi0957= 0;
    pi0958= 0;
    pi0959= 0;
    pi0960= 0;
    pi0961= 0;
    pi0962= 0;
    pi0963= 0;
    pi0964= 0;
    pi0965= 0;
    pi0966= 0;
    pi0967= 0;
    pi0968= 0;
    pi0969= 0;
    pi0970= 0;
    pi0971= 0;
    pi0972= 0;
    pi0973= 0;
    pi0974= 0;
    pi0975= 0;
    pi0976= 0;
    pi0977= 0;
    pi0978= 0;
    pi0979= 0;
    pi0980= 0;
    pi0981= 0;
    pi0982= 0;
    pi0983= 0;
    pi0984= 0;
    pi0985= 0;
    pi0986= 0;
    pi0987= 0;
    pi0988= 0;
    pi0989= 0;
    pi0990= 0;
    pi0991= 0;
    pi0992= 0;
    pi0993= 0;
    pi0994= 0;
    pi0995= 0;
    pi0996= 0;
    pi0997= 0;
    pi0998= 0;
    pi0999= 0;
    pi1000= 0;
    pi1001= 0;
    pi1002= 0;
    pi1003= 0;
    pi1004= 0;
    pi1005= 0;
    pi1006= 0;
    pi1007= 0;
    pi1008= 0;
    pi1009= 0;
    pi1010= 0;
    pi1011= 0;
    pi1012= 0;
    pi1013= 0;
    pi1014= 0;
    pi1015= 0;
    pi1016= 0;
    pi1017= 0;
    pi1018= 0;
    pi1019= 0;
    pi1020= 0;
    pi1021= 0;
    pi1022= 0;
    pi1023= 0;
    pi1024= 0;
    pi1025= 0;
    pi1026= 0;
    pi1027= 0;
    pi1028= 0;
    pi1029= 0;
    pi1030= 0;
    pi1031= 0;
    pi1032= 0;
    pi1033= 0;
    pi1034= 0;
    pi1035= 0;
    pi1036= 0;
    pi1037= 0;
    pi1038= 0;
    pi1039= 0;
    pi1040= 0;
    pi1041= 0;
    pi1042= 0;
    pi1043= 0;
    pi1044= 0;
    pi1045= 0;
    pi1046= 0;
    pi1047= 0;
    pi1048= 0;
    pi1049= 0;
    pi1050= 0;
    pi1051= 0;
    pi1052= 0;
    pi1053= 0;
    pi1054= 0;
    pi1055= 0;
    pi1056= 0;
    pi1057= 0;
    pi1058= 0;
    pi1059= 0;
    pi1060= 0;
    pi1061= 0;
    pi1062= 0;
    pi1063= 0;
    pi1064= 0;
    pi1065= 0;
    pi1066= 0;
    pi1067= 0;
    pi1068= 0;
    pi1069= 0;
    pi1070= 0;
    pi1071= 0;
    pi1072= 0;
    pi1073= 0;
    pi1074= 0;
    pi1075= 0;
    pi1076= 0;
    pi1077= 0;
    pi1078= 0;
    pi1079= 0;
    pi1080= 0;
    pi1081= 0;
    pi1082= 0;
    pi1083= 0;
    pi1084= 0;
    pi1085= 0;
    pi1086= 0;
    pi1087= 0;
    pi1088= 0;
    pi1089= 0;
    pi1090= 0;
    pi1091= 0;
    pi1092= 0;
    pi1093= 0;
    pi1094= 0;
    pi1095= 0;
    pi1096= 0;
    pi1097= 0;
    pi1098= 0;
    pi1099= 0;
    pi1100= 0;
    pi1101= 0;
    pi1102= 0;
    pi1103= 0;
    pi1104= 0;
    pi1105= 0;
    pi1106= 0;
    pi1107= 0;
    pi1108= 0;
    pi1109= 0;
    pi1110= 0;
    pi1111= 0;
    pi1112= 0;
    pi1113= 0;
    pi1114= 0;
    pi1115= 0;
    pi1116= 0;
    pi1117= 0;
    pi1118= 0;
    pi1119= 0;
    pi1120= 0;
    pi1121= 0;
    pi1122= 0;
    pi1123= 0;
    pi1124= 0;
    pi1125= 0;
    pi1126= 0;
    pi1127= 0;
    pi1128= 0;
    pi1129= 0;
    pi1130= 0;
    pi1131= 0;
    pi1132= 0;
    pi1133= 0;
    pi1134= 0;
    pi1135= 0;
    pi1136= 0;
    pi1137= 0;
    pi1138= 0;
    pi1139= 0;
    pi1140= 0;
    pi1141= 0;
    pi1142= 0;
    pi1143= 0;
    pi1144= 0;
    pi1145= 0;
    pi1146= 0;
    pi1147= 0;
    pi1148= 0;
    pi1149= 0;
    pi1150= 0;
    pi1151= 0;
    pi1152= 0;
    pi1153= 0;
    pi1154= 0;
    pi1155= 0;
    pi1156= 0;
    pi1157= 0;
    pi1158= 0;
    pi1159= 0;
    pi1160= 0;
    pi1161= 0;
    pi1162= 0;
    pi1163= 0;
    pi1164= 0;
    pi1165= 0;
    pi1166= 0;
    pi1167= 0;
    pi1168= 0;
    pi1169= 0;
    pi1170= 0;
    pi1171= 0;
    pi1172= 0;
    pi1173= 0;
    pi1174= 0;
    pi1175= 0;
    pi1176= 0;
    pi1177= 0;
    pi1178= 0;
    pi1179= 0;
    pi1180= 0;
    pi1181= 0;
    pi1182= 0;
    pi1183= 0;
    pi1184= 0;
    pi1185= 0;
    pi1186= 0;
    pi1187= 0;
    pi1188= 0;
    pi1189= 0;
    pi1190= 0;
    pi1191= 0;
    pi1192= 0;
    pi1193= 0;
    pi1194= 0;
    pi1195= 0;
    pi1196= 0;
    pi1197= 0;
    pi1198= 0;
    pi1199= 0;
    pi1200= 0;
    pi1201= 0;
    pi1202= 0;
    pi1203= 0;

    #10;

    for (i = 0; i < CYCLES; i = i + 1) begin
        // pi0000: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0000= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0000= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0000= (i + 0) % 2;  // Phase3: 翻转
          end
        end

        // pi0001: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0001= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0001= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0001= (i + 1) % 2;  // Phase3: 翻转
          end
        end

        // pi0002: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0002= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0002= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0002= (i + 2) % 2;  // Phase3: 翻转
          end
        end

        // pi0003: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0003= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0003= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0003= (i + 3) % 2;  // Phase3: 翻转
          end
        end

        // pi0004: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0004= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0004= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0004= (i + 4) % 2;  // Phase3: 翻转
          end
        end

        // pi0005: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0005= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0005= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0005= (i + 5) % 2;  // Phase3: 翻转
          end
        end

        // pi0006: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0006= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0006= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0006= (i + 6) % 2;  // Phase3: 翻转
          end
        end

        // pi0007: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0007= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0007= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0007= (i + 7) % 2;  // Phase3: 翻转
          end
        end

        // pi0008: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0008= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0008= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0008= (i + 8) % 2;  // Phase3: 翻转
          end
        end

        // pi0009: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0009= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0009= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0009= (i + 9) % 2;  // Phase3: 翻转
          end
        end

        // pi0010: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0010= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0010= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0010= (i + 10) % 2;  // Phase3: 翻转
          end
        end

        // pi0011: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0011= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0011= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0011= (i + 11) % 2;  // Phase3: 翻转
          end
        end

        // pi0012: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0012= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0012= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0012= (i + 12) % 2;  // Phase3: 翻转
          end
        end

        // pi0013: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0013= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0013= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0013= (i + 13) % 2;  // Phase3: 翻转
          end
        end

        // pi0014: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0014= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0014= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0014= (i + 14) % 2;  // Phase3: 翻转
          end
        end

        // pi0015: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0015= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0015= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0015= (i + 15) % 2;  // Phase3: 翻转
          end
        end

        // pi0016: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0016= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0016= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0016= (i + 16) % 2;  // Phase3: 翻转
          end
        end

        // pi0017: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0017= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0017= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0017= (i + 17) % 2;  // Phase3: 翻转
          end
        end

        // pi0018: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0018= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0018= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0018= (i + 18) % 2;  // Phase3: 翻转
          end
        end

        // pi0019: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0019= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0019= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0019= (i + 19) % 2;  // Phase3: 翻转
          end
        end

        // pi0020: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0020= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0020= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0020= (i + 20) % 2;  // Phase3: 翻转
          end
        end

        // pi0021: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0021= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0021= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0021= (i + 21) % 2;  // Phase3: 翻转
          end
        end

        // pi0022: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0022= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0022= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0022= (i + 22) % 2;  // Phase3: 翻转
          end
        end

        // pi0023: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0023= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0023= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0023= (i + 23) % 2;  // Phase3: 翻转
          end
        end

        // pi0024: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0024= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0024= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0024= (i + 24) % 2;  // Phase3: 翻转
          end
        end

        // pi0025: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0025= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0025= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0025= (i + 25) % 2;  // Phase3: 翻转
          end
        end

        // pi0026: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0026= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0026= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0026= (i + 26) % 2;  // Phase3: 翻转
          end
        end

        // pi0027: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0027= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0027= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0027= (i + 27) % 2;  // Phase3: 翻转
          end
        end

        // pi0028: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0028= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0028= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0028= (i + 28) % 2;  // Phase3: 翻转
          end
        end

        // pi0029: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0029= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0029= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0029= (i + 29) % 2;  // Phase3: 翻转
          end
        end

        // pi0030: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0030= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0030= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0030= (i + 30) % 2;  // Phase3: 翻转
          end
        end

        // pi0031: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0031= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0031= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0031= (i + 31) % 2;  // Phase3: 翻转
          end
        end

        // pi0032: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0032= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0032= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0032= (i + 32) % 2;  // Phase3: 翻转
          end
        end

        // pi0033: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0033= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0033= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0033= (i + 33) % 2;  // Phase3: 翻转
          end
        end

        // pi0034: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0034= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0034= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0034= (i + 34) % 2;  // Phase3: 翻转
          end
        end

        // pi0035: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0035= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0035= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0035= (i + 35) % 2;  // Phase3: 翻转
          end
        end

        // pi0036: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0036= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0036= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0036= (i + 36) % 2;  // Phase3: 翻转
          end
        end

        // pi0037: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0037= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0037= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0037= (i + 37) % 2;  // Phase3: 翻转
          end
        end

        // pi0038: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0038= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0038= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0038= (i + 38) % 2;  // Phase3: 翻转
          end
        end

        // pi0039: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0039= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0039= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0039= (i + 39) % 2;  // Phase3: 翻转
          end
        end

        // pi0040: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0040= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0040= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0040= (i + 40) % 2;  // Phase3: 翻转
          end
        end

        // pi0041: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0041= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0041= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0041= (i + 41) % 2;  // Phase3: 翻转
          end
        end

        // pi0042: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0042= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0042= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0042= (i + 42) % 2;  // Phase3: 翻转
          end
        end

        // pi0043: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0043= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0043= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0043= (i + 43) % 2;  // Phase3: 翻转
          end
        end

        // pi0044: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0044= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0044= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0044= (i + 44) % 2;  // Phase3: 翻转
          end
        end

        // pi0045: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0045= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0045= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0045= (i + 45) % 2;  // Phase3: 翻转
          end
        end

        // pi0046: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0046= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0046= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0046= (i + 46) % 2;  // Phase3: 翻转
          end
        end

        // pi0047: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0047= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0047= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0047= (i + 47) % 2;  // Phase3: 翻转
          end
        end

        // pi0048: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0048= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0048= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0048= (i + 48) % 2;  // Phase3: 翻转
          end
        end

        // pi0049: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0049= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0049= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0049= (i + 49) % 2;  // Phase3: 翻转
          end
        end

        // pi0050: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0050= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0050= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0050= (i + 50) % 2;  // Phase3: 翻转
          end
        end

        // pi0051: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0051= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0051= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0051= (i + 51) % 2;  // Phase3: 翻转
          end
        end

        // pi0052: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0052= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0052= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0052= (i + 52) % 2;  // Phase3: 翻转
          end
        end

        // pi0053: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0053= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0053= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0053= (i + 53) % 2;  // Phase3: 翻转
          end
        end

        // pi0054: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0054= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0054= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0054= (i + 54) % 2;  // Phase3: 翻转
          end
        end

        // pi0055: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0055= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0055= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0055= (i + 55) % 2;  // Phase3: 翻转
          end
        end

        // pi0056: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0056= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0056= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0056= (i + 56) % 2;  // Phase3: 翻转
          end
        end

        // pi0057: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0057= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0057= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0057= (i + 57) % 2;  // Phase3: 翻转
          end
        end

        // pi0058: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0058= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0058= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0058= (i + 58) % 2;  // Phase3: 翻转
          end
        end

        // pi0059: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0059= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0059= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0059= (i + 59) % 2;  // Phase3: 翻转
          end
        end

        // pi0060: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0060= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0060= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0060= (i + 60) % 2;  // Phase3: 翻转
          end
        end

        // pi0061: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0061= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0061= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0061= (i + 61) % 2;  // Phase3: 翻转
          end
        end

        // pi0062: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0062= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0062= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0062= (i + 62) % 2;  // Phase3: 翻转
          end
        end

        // pi0063: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0063= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0063= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0063= (i + 63) % 2;  // Phase3: 翻转
          end
        end

        // pi0064: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0064= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0064= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0064= (i + 64) % 2;  // Phase3: 翻转
          end
        end

        // pi0065: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0065= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0065= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0065= (i + 65) % 2;  // Phase3: 翻转
          end
        end

        // pi0066: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0066= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0066= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0066= (i + 66) % 2;  // Phase3: 翻转
          end
        end

        // pi0067: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0067= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0067= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0067= (i + 67) % 2;  // Phase3: 翻转
          end
        end

        // pi0068: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0068= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0068= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0068= (i + 68) % 2;  // Phase3: 翻转
          end
        end

        // pi0069: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0069= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0069= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0069= (i + 69) % 2;  // Phase3: 翻转
          end
        end

        // pi0070: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0070= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0070= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0070= (i + 70) % 2;  // Phase3: 翻转
          end
        end

        // pi0071: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0071= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0071= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0071= (i + 71) % 2;  // Phase3: 翻转
          end
        end

        // pi0072: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0072= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0072= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0072= (i + 72) % 2;  // Phase3: 翻转
          end
        end

        // pi0073: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0073= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0073= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0073= (i + 73) % 2;  // Phase3: 翻转
          end
        end

        // pi0074: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0074= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0074= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0074= (i + 74) % 2;  // Phase3: 翻转
          end
        end

        // pi0075: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0075= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0075= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0075= (i + 75) % 2;  // Phase3: 翻转
          end
        end

        // pi0076: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0076= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0076= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0076= (i + 76) % 2;  // Phase3: 翻转
          end
        end

        // pi0077: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0077= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0077= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0077= (i + 77) % 2;  // Phase3: 翻转
          end
        end

        // pi0078: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0078= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0078= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0078= (i + 78) % 2;  // Phase3: 翻转
          end
        end

        // pi0079: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0079= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0079= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0079= (i + 79) % 2;  // Phase3: 翻转
          end
        end

        // pi0080: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0080= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0080= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0080= (i + 80) % 2;  // Phase3: 翻转
          end
        end

        // pi0081: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0081= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0081= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0081= (i + 81) % 2;  // Phase3: 翻转
          end
        end

        // pi0082: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0082= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0082= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0082= (i + 82) % 2;  // Phase3: 翻转
          end
        end

        // pi0083: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0083= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0083= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0083= (i + 83) % 2;  // Phase3: 翻转
          end
        end

        // pi0084: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0084= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0084= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0084= (i + 84) % 2;  // Phase3: 翻转
          end
        end

        // pi0085: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0085= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0085= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0085= (i + 85) % 2;  // Phase3: 翻转
          end
        end

        // pi0086: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0086= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0086= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0086= (i + 86) % 2;  // Phase3: 翻转
          end
        end

        // pi0087: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0087= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0087= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0087= (i + 87) % 2;  // Phase3: 翻转
          end
        end

        // pi0088: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0088= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0088= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0088= (i + 88) % 2;  // Phase3: 翻转
          end
        end

        // pi0089: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0089= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0089= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0089= (i + 89) % 2;  // Phase3: 翻转
          end
        end

        // pi0090: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0090= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0090= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0090= (i + 90) % 2;  // Phase3: 翻转
          end
        end

        // pi0091: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0091= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0091= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0091= (i + 91) % 2;  // Phase3: 翻转
          end
        end

        // pi0092: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0092= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0092= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0092= (i + 92) % 2;  // Phase3: 翻转
          end
        end

        // pi0093: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0093= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0093= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0093= (i + 93) % 2;  // Phase3: 翻转
          end
        end

        // pi0094: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0094= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0094= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0094= (i + 94) % 2;  // Phase3: 翻转
          end
        end

        // pi0095: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0095= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0095= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0095= (i + 95) % 2;  // Phase3: 翻转
          end
        end

        // pi0096: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0096= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0096= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0096= (i + 96) % 2;  // Phase3: 翻转
          end
        end

        // pi0097: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0097= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0097= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0097= (i + 97) % 2;  // Phase3: 翻转
          end
        end

        // pi0098: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0098= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0098= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0098= (i + 98) % 2;  // Phase3: 翻转
          end
        end

        // pi0099: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0099= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0099= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0099= (i + 99) % 2;  // Phase3: 翻转
          end
        end

        // pi0100: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0100= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0100= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0100= (i + 100) % 2;  // Phase3: 翻转
          end
        end

        // pi0101: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0101= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0101= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0101= (i + 101) % 2;  // Phase3: 翻转
          end
        end

        // pi0102: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0102= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0102= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0102= (i + 102) % 2;  // Phase3: 翻转
          end
        end

        // pi0103: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0103= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0103= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0103= (i + 103) % 2;  // Phase3: 翻转
          end
        end

        // pi0104: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0104= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0104= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0104= (i + 104) % 2;  // Phase3: 翻转
          end
        end

        // pi0105: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0105= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0105= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0105= (i + 105) % 2;  // Phase3: 翻转
          end
        end

        // pi0106: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0106= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0106= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0106= (i + 106) % 2;  // Phase3: 翻转
          end
        end

        // pi0107: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0107= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0107= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0107= (i + 107) % 2;  // Phase3: 翻转
          end
        end

        // pi0108: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0108= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0108= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0108= (i + 108) % 2;  // Phase3: 翻转
          end
        end

        // pi0109: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0109= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0109= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0109= (i + 109) % 2;  // Phase3: 翻转
          end
        end

        // pi0110: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0110= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0110= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0110= (i + 110) % 2;  // Phase3: 翻转
          end
        end

        // pi0111: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0111= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0111= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0111= (i + 111) % 2;  // Phase3: 翻转
          end
        end

        // pi0112: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0112= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0112= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0112= (i + 112) % 2;  // Phase3: 翻转
          end
        end

        // pi0113: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0113= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0113= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0113= (i + 113) % 2;  // Phase3: 翻转
          end
        end

        // pi0114: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0114= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0114= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0114= (i + 114) % 2;  // Phase3: 翻转
          end
        end

        // pi0115: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0115= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0115= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0115= (i + 115) % 2;  // Phase3: 翻转
          end
        end

        // pi0116: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0116= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0116= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0116= (i + 116) % 2;  // Phase3: 翻转
          end
        end

        // pi0117: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0117= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0117= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0117= (i + 117) % 2;  // Phase3: 翻转
          end
        end

        // pi0118: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0118= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0118= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0118= (i + 118) % 2;  // Phase3: 翻转
          end
        end

        // pi0119: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0119= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0119= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0119= (i + 119) % 2;  // Phase3: 翻转
          end
        end

        // pi0120: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0120= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0120= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0120= (i + 120) % 2;  // Phase3: 翻转
          end
        end

        // pi0121: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0121= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0121= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0121= (i + 121) % 2;  // Phase3: 翻转
          end
        end

        // pi0122: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0122= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0122= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0122= (i + 122) % 2;  // Phase3: 翻转
          end
        end

        // pi0123: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0123= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0123= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0123= (i + 123) % 2;  // Phase3: 翻转
          end
        end

        // pi0124: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0124= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0124= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0124= (i + 124) % 2;  // Phase3: 翻转
          end
        end

        // pi0125: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0125= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0125= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0125= (i + 125) % 2;  // Phase3: 翻转
          end
        end

        // pi0126: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0126= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0126= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0126= (i + 126) % 2;  // Phase3: 翻转
          end
        end

        // pi0127: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0127= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0127= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0127= (i + 127) % 2;  // Phase3: 翻转
          end
        end

        // pi0128: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0128= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0128= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0128= (i + 128) % 2;  // Phase3: 翻转
          end
        end

        // pi0129: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0129= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0129= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0129= (i + 129) % 2;  // Phase3: 翻转
          end
        end

        // pi0130: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0130= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0130= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0130= (i + 130) % 2;  // Phase3: 翻转
          end
        end

        // pi0131: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0131= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0131= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0131= (i + 131) % 2;  // Phase3: 翻转
          end
        end

        // pi0132: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0132= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0132= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0132= (i + 132) % 2;  // Phase3: 翻转
          end
        end

        // pi0133: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0133= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0133= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0133= (i + 133) % 2;  // Phase3: 翻转
          end
        end

        // pi0134: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0134= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0134= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0134= (i + 134) % 2;  // Phase3: 翻转
          end
        end

        // pi0135: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0135= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0135= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0135= (i + 135) % 2;  // Phase3: 翻转
          end
        end

        // pi0136: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0136= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0136= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0136= (i + 136) % 2;  // Phase3: 翻转
          end
        end

        // pi0137: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0137= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0137= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0137= (i + 137) % 2;  // Phase3: 翻转
          end
        end

        // pi0138: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0138= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0138= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0138= (i + 138) % 2;  // Phase3: 翻转
          end
        end

        // pi0139: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0139= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0139= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0139= (i + 139) % 2;  // Phase3: 翻转
          end
        end

        // pi0140: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0140= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0140= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0140= (i + 140) % 2;  // Phase3: 翻转
          end
        end

        // pi0141: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0141= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0141= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0141= (i + 141) % 2;  // Phase3: 翻转
          end
        end

        // pi0142: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0142= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0142= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0142= (i + 142) % 2;  // Phase3: 翻转
          end
        end

        // pi0143: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0143= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0143= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0143= (i + 143) % 2;  // Phase3: 翻转
          end
        end

        // pi0144: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0144= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0144= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0144= (i + 144) % 2;  // Phase3: 翻转
          end
        end

        // pi0145: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0145= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0145= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0145= (i + 145) % 2;  // Phase3: 翻转
          end
        end

        // pi0146: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0146= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0146= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0146= (i + 146) % 2;  // Phase3: 翻转
          end
        end

        // pi0147: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0147= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0147= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0147= (i + 147) % 2;  // Phase3: 翻转
          end
        end

        // pi0148: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0148= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0148= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0148= (i + 148) % 2;  // Phase3: 翻转
          end
        end

        // pi0149: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0149= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0149= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0149= (i + 149) % 2;  // Phase3: 翻转
          end
        end

        // pi0150: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0150= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0150= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0150= (i + 150) % 2;  // Phase3: 翻转
          end
        end

        // pi0151: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0151= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0151= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0151= (i + 151) % 2;  // Phase3: 翻转
          end
        end

        // pi0152: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0152= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0152= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0152= (i + 152) % 2;  // Phase3: 翻转
          end
        end

        // pi0153: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0153= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0153= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0153= (i + 153) % 2;  // Phase3: 翻转
          end
        end

        // pi0154: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0154= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0154= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0154= (i + 154) % 2;  // Phase3: 翻转
          end
        end

        // pi0155: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0155= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0155= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0155= (i + 155) % 2;  // Phase3: 翻转
          end
        end

        // pi0156: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0156= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0156= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0156= (i + 156) % 2;  // Phase3: 翻转
          end
        end

        // pi0157: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0157= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0157= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0157= (i + 157) % 2;  // Phase3: 翻转
          end
        end

        // pi0158: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0158= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0158= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0158= (i + 158) % 2;  // Phase3: 翻转
          end
        end

        // pi0159: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0159= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0159= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0159= (i + 159) % 2;  // Phase3: 翻转
          end
        end

        // pi0160: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0160= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0160= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0160= (i + 160) % 2;  // Phase3: 翻转
          end
        end

        // pi0161: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0161= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0161= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0161= (i + 161) % 2;  // Phase3: 翻转
          end
        end

        // pi0162: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0162= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0162= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0162= (i + 162) % 2;  // Phase3: 翻转
          end
        end

        // pi0163: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0163= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0163= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0163= (i + 163) % 2;  // Phase3: 翻转
          end
        end

        // pi0164: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0164= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0164= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0164= (i + 164) % 2;  // Phase3: 翻转
          end
        end

        // pi0165: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0165= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0165= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0165= (i + 165) % 2;  // Phase3: 翻转
          end
        end

        // pi0166: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0166= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0166= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0166= (i + 166) % 2;  // Phase3: 翻转
          end
        end

        // pi0167: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0167= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0167= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0167= (i + 167) % 2;  // Phase3: 翻转
          end
        end

        // pi0168: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0168= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0168= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0168= (i + 168) % 2;  // Phase3: 翻转
          end
        end

        // pi0169: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0169= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0169= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0169= (i + 169) % 2;  // Phase3: 翻转
          end
        end

        // pi0170: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0170= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0170= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0170= (i + 170) % 2;  // Phase3: 翻转
          end
        end

        // pi0171: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0171= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0171= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0171= (i + 171) % 2;  // Phase3: 翻转
          end
        end

        // pi0172: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0172= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0172= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0172= (i + 172) % 2;  // Phase3: 翻转
          end
        end

        // pi0173: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0173= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0173= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0173= (i + 173) % 2;  // Phase3: 翻转
          end
        end

        // pi0174: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0174= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0174= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0174= (i + 174) % 2;  // Phase3: 翻转
          end
        end

        // pi0175: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0175= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0175= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0175= (i + 175) % 2;  // Phase3: 翻转
          end
        end

        // pi0176: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0176= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0176= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0176= (i + 176) % 2;  // Phase3: 翻转
          end
        end

        // pi0177: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0177= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0177= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0177= (i + 177) % 2;  // Phase3: 翻转
          end
        end

        // pi0178: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0178= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0178= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0178= (i + 178) % 2;  // Phase3: 翻转
          end
        end

        // pi0179: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0179= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0179= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0179= (i + 179) % 2;  // Phase3: 翻转
          end
        end

        // pi0180: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0180= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0180= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0180= (i + 180) % 2;  // Phase3: 翻转
          end
        end

        // pi0181: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0181= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0181= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0181= (i + 181) % 2;  // Phase3: 翻转
          end
        end

        // pi0182: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0182= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0182= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0182= (i + 182) % 2;  // Phase3: 翻转
          end
        end

        // pi0183: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0183= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0183= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0183= (i + 183) % 2;  // Phase3: 翻转
          end
        end

        // pi0184: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0184= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0184= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0184= (i + 184) % 2;  // Phase3: 翻转
          end
        end

        // pi0185: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0185= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0185= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0185= (i + 185) % 2;  // Phase3: 翻转
          end
        end

        // pi0186: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0186= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0186= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0186= (i + 186) % 2;  // Phase3: 翻转
          end
        end

        // pi0187: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0187= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0187= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0187= (i + 187) % 2;  // Phase3: 翻转
          end
        end

        // pi0188: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0188= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0188= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0188= (i + 188) % 2;  // Phase3: 翻转
          end
        end

        // pi0189: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0189= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0189= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0189= (i + 189) % 2;  // Phase3: 翻转
          end
        end

        // pi0190: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0190= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0190= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0190= (i + 190) % 2;  // Phase3: 翻转
          end
        end

        // pi0191: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0191= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0191= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0191= (i + 191) % 2;  // Phase3: 翻转
          end
        end

        // pi0192: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0192= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0192= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0192= (i + 192) % 2;  // Phase3: 翻转
          end
        end

        // pi0193: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0193= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0193= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0193= (i + 193) % 2;  // Phase3: 翻转
          end
        end

        // pi0194: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0194= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0194= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0194= (i + 194) % 2;  // Phase3: 翻转
          end
        end

        // pi0195: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0195= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0195= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0195= (i + 195) % 2;  // Phase3: 翻转
          end
        end

        // pi0196: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0196= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0196= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0196= (i + 196) % 2;  // Phase3: 翻转
          end
        end

        // pi0197: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0197= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0197= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0197= (i + 197) % 2;  // Phase3: 翻转
          end
        end

        // pi0198: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0198= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0198= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0198= (i + 198) % 2;  // Phase3: 翻转
          end
        end

        // pi0199: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0199= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0199= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0199= (i + 199) % 2;  // Phase3: 翻转
          end
        end

        // pi0200: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0200= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0200= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0200= (i + 200) % 2;  // Phase3: 翻转
          end
        end

        // pi0201: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0201= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0201= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0201= (i + 201) % 2;  // Phase3: 翻转
          end
        end

        // pi0202: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0202= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0202= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0202= (i + 202) % 2;  // Phase3: 翻转
          end
        end

        // pi0203: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0203= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0203= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0203= (i + 203) % 2;  // Phase3: 翻转
          end
        end

        // pi0204: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0204= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0204= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0204= (i + 204) % 2;  // Phase3: 翻转
          end
        end

        // pi0205: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0205= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0205= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0205= (i + 205) % 2;  // Phase3: 翻转
          end
        end

        // pi0206: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0206= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0206= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0206= (i + 206) % 2;  // Phase3: 翻转
          end
        end

        // pi0207: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0207= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0207= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0207= (i + 207) % 2;  // Phase3: 翻转
          end
        end

        // pi0208: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0208= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0208= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0208= (i + 208) % 2;  // Phase3: 翻转
          end
        end

        // pi0209: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0209= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0209= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0209= (i + 209) % 2;  // Phase3: 翻转
          end
        end

        // pi0210: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0210= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0210= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0210= (i + 210) % 2;  // Phase3: 翻转
          end
        end

        // pi0211: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0211= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0211= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0211= (i + 211) % 2;  // Phase3: 翻转
          end
        end

        // pi0212: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0212= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0212= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0212= (i + 212) % 2;  // Phase3: 翻转
          end
        end

        // pi0213: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0213= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0213= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0213= (i + 213) % 2;  // Phase3: 翻转
          end
        end

        // pi0214: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0214= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0214= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0214= (i + 214) % 2;  // Phase3: 翻转
          end
        end

        // pi0215: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0215= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0215= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0215= (i + 215) % 2;  // Phase3: 翻转
          end
        end

        // pi0216: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0216= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0216= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0216= (i + 216) % 2;  // Phase3: 翻转
          end
        end

        // pi0217: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0217= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0217= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0217= (i + 217) % 2;  // Phase3: 翻转
          end
        end

        // pi0218: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0218= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0218= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0218= (i + 218) % 2;  // Phase3: 翻转
          end
        end

        // pi0219: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0219= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0219= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0219= (i + 219) % 2;  // Phase3: 翻转
          end
        end

        // pi0220: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0220= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0220= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0220= (i + 220) % 2;  // Phase3: 翻转
          end
        end

        // pi0221: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0221= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0221= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0221= (i + 221) % 2;  // Phase3: 翻转
          end
        end

        // pi0222: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0222= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0222= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0222= (i + 222) % 2;  // Phase3: 翻转
          end
        end

        // pi0223: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0223= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0223= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0223= (i + 223) % 2;  // Phase3: 翻转
          end
        end

        // pi0224: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0224= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0224= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0224= (i + 224) % 2;  // Phase3: 翻转
          end
        end

        // pi0225: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0225= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0225= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0225= (i + 225) % 2;  // Phase3: 翻转
          end
        end

        // pi0226: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0226= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0226= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0226= (i + 226) % 2;  // Phase3: 翻转
          end
        end

        // pi0227: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0227= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0227= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0227= (i + 227) % 2;  // Phase3: 翻转
          end
        end

        // pi0228: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0228= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0228= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0228= (i + 228) % 2;  // Phase3: 翻转
          end
        end

        // pi0229: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0229= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0229= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0229= (i + 229) % 2;  // Phase3: 翻转
          end
        end

        // pi0230: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0230= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0230= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0230= (i + 230) % 2;  // Phase3: 翻转
          end
        end

        // pi0231: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0231= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0231= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0231= (i + 231) % 2;  // Phase3: 翻转
          end
        end

        // pi0232: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0232= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0232= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0232= (i + 232) % 2;  // Phase3: 翻转
          end
        end

        // pi0233: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0233= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0233= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0233= (i + 233) % 2;  // Phase3: 翻转
          end
        end

        // pi0234: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0234= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0234= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0234= (i + 234) % 2;  // Phase3: 翻转
          end
        end

        // pi0235: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0235= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0235= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0235= (i + 235) % 2;  // Phase3: 翻转
          end
        end

        // pi0236: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0236= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0236= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0236= (i + 236) % 2;  // Phase3: 翻转
          end
        end

        // pi0237: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0237= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0237= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0237= (i + 237) % 2;  // Phase3: 翻转
          end
        end

        // pi0238: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0238= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0238= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0238= (i + 238) % 2;  // Phase3: 翻转
          end
        end

        // pi0239: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0239= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0239= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0239= (i + 239) % 2;  // Phase3: 翻转
          end
        end

        // pi0240: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0240= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0240= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0240= (i + 240) % 2;  // Phase3: 翻转
          end
        end

        // pi0241: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0241= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0241= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0241= (i + 241) % 2;  // Phase3: 翻转
          end
        end

        // pi0242: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0242= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0242= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0242= (i + 242) % 2;  // Phase3: 翻转
          end
        end

        // pi0243: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0243= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0243= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0243= (i + 243) % 2;  // Phase3: 翻转
          end
        end

        // pi0244: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0244= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0244= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0244= (i + 244) % 2;  // Phase3: 翻转
          end
        end

        // pi0245: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0245= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0245= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0245= (i + 245) % 2;  // Phase3: 翻转
          end
        end

        // pi0246: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0246= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0246= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0246= (i + 246) % 2;  // Phase3: 翻转
          end
        end

        // pi0247: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0247= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0247= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0247= (i + 247) % 2;  // Phase3: 翻转
          end
        end

        // pi0248: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0248= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0248= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0248= (i + 248) % 2;  // Phase3: 翻转
          end
        end

        // pi0249: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0249= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0249= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0249= (i + 249) % 2;  // Phase3: 翻转
          end
        end

        // pi0250: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0250= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0250= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0250= (i + 250) % 2;  // Phase3: 翻转
          end
        end

        // pi0251: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0251= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0251= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0251= (i + 251) % 2;  // Phase3: 翻转
          end
        end

        // pi0252: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0252= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0252= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0252= (i + 252) % 2;  // Phase3: 翻转
          end
        end

        // pi0253: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0253= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0253= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0253= (i + 253) % 2;  // Phase3: 翻转
          end
        end

        // pi0254: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0254= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0254= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0254= (i + 254) % 2;  // Phase3: 翻转
          end
        end

        // pi0255: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0255= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0255= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0255= (i + 255) % 2;  // Phase3: 翻转
          end
        end

        // pi0256: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0256= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0256= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0256= (i + 256) % 2;  // Phase3: 翻转
          end
        end

        // pi0257: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0257= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0257= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0257= (i + 257) % 2;  // Phase3: 翻转
          end
        end

        // pi0258: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0258= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0258= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0258= (i + 258) % 2;  // Phase3: 翻转
          end
        end

        // pi0259: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0259= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0259= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0259= (i + 259) % 2;  // Phase3: 翻转
          end
        end

        // pi0260: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0260= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0260= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0260= (i + 260) % 2;  // Phase3: 翻转
          end
        end

        // pi0261: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0261= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0261= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0261= (i + 261) % 2;  // Phase3: 翻转
          end
        end

        // pi0262: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0262= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0262= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0262= (i + 262) % 2;  // Phase3: 翻转
          end
        end

        // pi0263: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0263= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0263= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0263= (i + 263) % 2;  // Phase3: 翻转
          end
        end

        // pi0264: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0264= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0264= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0264= (i + 264) % 2;  // Phase3: 翻转
          end
        end

        // pi0265: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0265= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0265= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0265= (i + 265) % 2;  // Phase3: 翻转
          end
        end

        // pi0266: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0266= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0266= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0266= (i + 266) % 2;  // Phase3: 翻转
          end
        end

        // pi0267: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0267= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0267= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0267= (i + 267) % 2;  // Phase3: 翻转
          end
        end

        // pi0268: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0268= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0268= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0268= (i + 268) % 2;  // Phase3: 翻转
          end
        end

        // pi0269: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0269= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0269= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0269= (i + 269) % 2;  // Phase3: 翻转
          end
        end

        // pi0270: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0270= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0270= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0270= (i + 270) % 2;  // Phase3: 翻转
          end
        end

        // pi0271: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0271= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0271= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0271= (i + 271) % 2;  // Phase3: 翻转
          end
        end

        // pi0272: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0272= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0272= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0272= (i + 272) % 2;  // Phase3: 翻转
          end
        end

        // pi0273: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0273= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0273= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0273= (i + 273) % 2;  // Phase3: 翻转
          end
        end

        // pi0274: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0274= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0274= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0274= (i + 274) % 2;  // Phase3: 翻转
          end
        end

        // pi0275: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0275= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0275= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0275= (i + 275) % 2;  // Phase3: 翻转
          end
        end

        // pi0276: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0276= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0276= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0276= (i + 276) % 2;  // Phase3: 翻转
          end
        end

        // pi0277: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0277= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0277= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0277= (i + 277) % 2;  // Phase3: 翻转
          end
        end

        // pi0278: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0278= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0278= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0278= (i + 278) % 2;  // Phase3: 翻转
          end
        end

        // pi0279: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0279= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0279= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0279= (i + 279) % 2;  // Phase3: 翻转
          end
        end

        // pi0280: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0280= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0280= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0280= (i + 280) % 2;  // Phase3: 翻转
          end
        end

        // pi0281: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0281= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0281= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0281= (i + 281) % 2;  // Phase3: 翻转
          end
        end

        // pi0282: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0282= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0282= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0282= (i + 282) % 2;  // Phase3: 翻转
          end
        end

        // pi0283: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0283= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0283= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0283= (i + 283) % 2;  // Phase3: 翻转
          end
        end

        // pi0284: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0284= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0284= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0284= (i + 284) % 2;  // Phase3: 翻转
          end
        end

        // pi0285: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0285= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0285= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0285= (i + 285) % 2;  // Phase3: 翻转
          end
        end

        // pi0286: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0286= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0286= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0286= (i + 286) % 2;  // Phase3: 翻转
          end
        end

        // pi0287: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0287= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0287= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0287= (i + 287) % 2;  // Phase3: 翻转
          end
        end

        // pi0288: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0288= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0288= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0288= (i + 288) % 2;  // Phase3: 翻转
          end
        end

        // pi0289: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0289= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0289= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0289= (i + 289) % 2;  // Phase3: 翻转
          end
        end

        // pi0290: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0290= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0290= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0290= (i + 290) % 2;  // Phase3: 翻转
          end
        end

        // pi0291: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0291= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0291= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0291= (i + 291) % 2;  // Phase3: 翻转
          end
        end

        // pi0292: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0292= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0292= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0292= (i + 292) % 2;  // Phase3: 翻转
          end
        end

        // pi0293: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0293= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0293= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0293= (i + 293) % 2;  // Phase3: 翻转
          end
        end

        // pi0294: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0294= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0294= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0294= (i + 294) % 2;  // Phase3: 翻转
          end
        end

        // pi0295: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0295= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0295= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0295= (i + 295) % 2;  // Phase3: 翻转
          end
        end

        // pi0296: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0296= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0296= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0296= (i + 296) % 2;  // Phase3: 翻转
          end
        end

        // pi0297: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0297= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0297= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0297= (i + 297) % 2;  // Phase3: 翻转
          end
        end

        // pi0298: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0298= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0298= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0298= (i + 298) % 2;  // Phase3: 翻转
          end
        end

        // pi0299: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0299= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0299= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0299= (i + 299) % 2;  // Phase3: 翻转
          end
        end

        // pi0300: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0300= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0300= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0300= (i + 300) % 2;  // Phase3: 翻转
          end
        end

        // pi0301: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0301= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0301= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0301= (i + 301) % 2;  // Phase3: 翻转
          end
        end

        // pi0302: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0302= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0302= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0302= (i + 302) % 2;  // Phase3: 翻转
          end
        end

        // pi0303: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0303= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0303= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0303= (i + 303) % 2;  // Phase3: 翻转
          end
        end

        // pi0304: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0304= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0304= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0304= (i + 304) % 2;  // Phase3: 翻转
          end
        end

        // pi0305: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0305= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0305= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0305= (i + 305) % 2;  // Phase3: 翻转
          end
        end

        // pi0306: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0306= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0306= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0306= (i + 306) % 2;  // Phase3: 翻转
          end
        end

        // pi0307: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0307= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0307= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0307= (i + 307) % 2;  // Phase3: 翻转
          end
        end

        // pi0308: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0308= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0308= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0308= (i + 308) % 2;  // Phase3: 翻转
          end
        end

        // pi0309: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0309= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0309= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0309= (i + 309) % 2;  // Phase3: 翻转
          end
        end

        // pi0310: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0310= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0310= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0310= (i + 310) % 2;  // Phase3: 翻转
          end
        end

        // pi0311: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0311= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0311= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0311= (i + 311) % 2;  // Phase3: 翻转
          end
        end

        // pi0312: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0312= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0312= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0312= (i + 312) % 2;  // Phase3: 翻转
          end
        end

        // pi0313: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0313= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0313= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0313= (i + 313) % 2;  // Phase3: 翻转
          end
        end

        // pi0314: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0314= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0314= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0314= (i + 314) % 2;  // Phase3: 翻转
          end
        end

        // pi0315: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0315= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0315= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0315= (i + 315) % 2;  // Phase3: 翻转
          end
        end

        // pi0316: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0316= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0316= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0316= (i + 316) % 2;  // Phase3: 翻转
          end
        end

        // pi0317: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0317= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0317= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0317= (i + 317) % 2;  // Phase3: 翻转
          end
        end

        // pi0318: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0318= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0318= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0318= (i + 318) % 2;  // Phase3: 翻转
          end
        end

        // pi0319: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0319= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0319= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0319= (i + 319) % 2;  // Phase3: 翻转
          end
        end

        // pi0320: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0320= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0320= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0320= (i + 320) % 2;  // Phase3: 翻转
          end
        end

        // pi0321: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0321= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0321= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0321= (i + 321) % 2;  // Phase3: 翻转
          end
        end

        // pi0322: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0322= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0322= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0322= (i + 322) % 2;  // Phase3: 翻转
          end
        end

        // pi0323: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0323= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0323= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0323= (i + 323) % 2;  // Phase3: 翻转
          end
        end

        // pi0324: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0324= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0324= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0324= (i + 324) % 2;  // Phase3: 翻转
          end
        end

        // pi0325: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0325= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0325= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0325= (i + 325) % 2;  // Phase3: 翻转
          end
        end

        // pi0326: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0326= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0326= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0326= (i + 326) % 2;  // Phase3: 翻转
          end
        end

        // pi0327: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0327= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0327= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0327= (i + 327) % 2;  // Phase3: 翻转
          end
        end

        // pi0328: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0328= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0328= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0328= (i + 328) % 2;  // Phase3: 翻转
          end
        end

        // pi0329: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0329= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0329= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0329= (i + 329) % 2;  // Phase3: 翻转
          end
        end

        // pi0330: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0330= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0330= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0330= (i + 330) % 2;  // Phase3: 翻转
          end
        end

        // pi0331: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0331= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0331= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0331= (i + 331) % 2;  // Phase3: 翻转
          end
        end

        // pi0332: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0332= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0332= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0332= (i + 332) % 2;  // Phase3: 翻转
          end
        end

        // pi0333: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0333= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0333= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0333= (i + 333) % 2;  // Phase3: 翻转
          end
        end

        // pi0334: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0334= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0334= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0334= (i + 334) % 2;  // Phase3: 翻转
          end
        end

        // pi0335: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0335= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0335= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0335= (i + 335) % 2;  // Phase3: 翻转
          end
        end

        // pi0336: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0336= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0336= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0336= (i + 336) % 2;  // Phase3: 翻转
          end
        end

        // pi0337: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0337= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0337= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0337= (i + 337) % 2;  // Phase3: 翻转
          end
        end

        // pi0338: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0338= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0338= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0338= (i + 338) % 2;  // Phase3: 翻转
          end
        end

        // pi0339: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0339= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0339= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0339= (i + 339) % 2;  // Phase3: 翻转
          end
        end

        // pi0340: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0340= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0340= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0340= (i + 340) % 2;  // Phase3: 翻转
          end
        end

        // pi0341: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0341= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0341= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0341= (i + 341) % 2;  // Phase3: 翻转
          end
        end

        // pi0342: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0342= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0342= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0342= (i + 342) % 2;  // Phase3: 翻转
          end
        end

        // pi0343: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0343= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0343= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0343= (i + 343) % 2;  // Phase3: 翻转
          end
        end

        // pi0344: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0344= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0344= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0344= (i + 344) % 2;  // Phase3: 翻转
          end
        end

        // pi0345: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0345= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0345= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0345= (i + 345) % 2;  // Phase3: 翻转
          end
        end

        // pi0346: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0346= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0346= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0346= (i + 346) % 2;  // Phase3: 翻转
          end
        end

        // pi0347: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0347= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0347= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0347= (i + 347) % 2;  // Phase3: 翻转
          end
        end

        // pi0348: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0348= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0348= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0348= (i + 348) % 2;  // Phase3: 翻转
          end
        end

        // pi0349: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0349= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0349= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0349= (i + 349) % 2;  // Phase3: 翻转
          end
        end

        // pi0350: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0350= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0350= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0350= (i + 350) % 2;  // Phase3: 翻转
          end
        end

        // pi0351: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0351= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0351= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0351= (i + 351) % 2;  // Phase3: 翻转
          end
        end

        // pi0352: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0352= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0352= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0352= (i + 352) % 2;  // Phase3: 翻转
          end
        end

        // pi0353: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0353= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0353= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0353= (i + 353) % 2;  // Phase3: 翻转
          end
        end

        // pi0354: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0354= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0354= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0354= (i + 354) % 2;  // Phase3: 翻转
          end
        end

        // pi0355: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0355= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0355= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0355= (i + 355) % 2;  // Phase3: 翻转
          end
        end

        // pi0356: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0356= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0356= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0356= (i + 356) % 2;  // Phase3: 翻转
          end
        end

        // pi0357: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0357= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0357= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0357= (i + 357) % 2;  // Phase3: 翻转
          end
        end

        // pi0358: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0358= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0358= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0358= (i + 358) % 2;  // Phase3: 翻转
          end
        end

        // pi0359: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0359= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0359= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0359= (i + 359) % 2;  // Phase3: 翻转
          end
        end

        // pi0360: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0360= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0360= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0360= (i + 360) % 2;  // Phase3: 翻转
          end
        end

        // pi0361: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0361= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0361= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0361= (i + 361) % 2;  // Phase3: 翻转
          end
        end

        // pi0362: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0362= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0362= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0362= (i + 362) % 2;  // Phase3: 翻转
          end
        end

        // pi0363: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0363= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0363= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0363= (i + 363) % 2;  // Phase3: 翻转
          end
        end

        // pi0364: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0364= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0364= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0364= (i + 364) % 2;  // Phase3: 翻转
          end
        end

        // pi0365: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0365= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0365= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0365= (i + 365) % 2;  // Phase3: 翻转
          end
        end

        // pi0366: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0366= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0366= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0366= (i + 366) % 2;  // Phase3: 翻转
          end
        end

        // pi0367: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0367= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0367= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0367= (i + 367) % 2;  // Phase3: 翻转
          end
        end

        // pi0368: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0368= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0368= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0368= (i + 368) % 2;  // Phase3: 翻转
          end
        end

        // pi0369: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0369= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0369= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0369= (i + 369) % 2;  // Phase3: 翻转
          end
        end

        // pi0370: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0370= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0370= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0370= (i + 370) % 2;  // Phase3: 翻转
          end
        end

        // pi0371: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0371= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0371= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0371= (i + 371) % 2;  // Phase3: 翻转
          end
        end

        // pi0372: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0372= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0372= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0372= (i + 372) % 2;  // Phase3: 翻转
          end
        end

        // pi0373: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0373= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0373= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0373= (i + 373) % 2;  // Phase3: 翻转
          end
        end

        // pi0374: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0374= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0374= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0374= (i + 374) % 2;  // Phase3: 翻转
          end
        end

        // pi0375: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0375= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0375= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0375= (i + 375) % 2;  // Phase3: 翻转
          end
        end

        // pi0376: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0376= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0376= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0376= (i + 376) % 2;  // Phase3: 翻转
          end
        end

        // pi0377: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0377= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0377= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0377= (i + 377) % 2;  // Phase3: 翻转
          end
        end

        // pi0378: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0378= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0378= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0378= (i + 378) % 2;  // Phase3: 翻转
          end
        end

        // pi0379: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0379= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0379= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0379= (i + 379) % 2;  // Phase3: 翻转
          end
        end

        // pi0380: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0380= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0380= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0380= (i + 380) % 2;  // Phase3: 翻转
          end
        end

        // pi0381: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0381= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0381= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0381= (i + 381) % 2;  // Phase3: 翻转
          end
        end

        // pi0382: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0382= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0382= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0382= (i + 382) % 2;  // Phase3: 翻转
          end
        end

        // pi0383: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0383= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0383= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0383= (i + 383) % 2;  // Phase3: 翻转
          end
        end

        // pi0384: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0384= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0384= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0384= (i + 384) % 2;  // Phase3: 翻转
          end
        end

        // pi0385: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0385= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0385= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0385= (i + 385) % 2;  // Phase3: 翻转
          end
        end

        // pi0386: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0386= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0386= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0386= (i + 386) % 2;  // Phase3: 翻转
          end
        end

        // pi0387: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0387= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0387= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0387= (i + 387) % 2;  // Phase3: 翻转
          end
        end

        // pi0388: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0388= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0388= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0388= (i + 388) % 2;  // Phase3: 翻转
          end
        end

        // pi0389: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0389= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0389= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0389= (i + 389) % 2;  // Phase3: 翻转
          end
        end

        // pi0390: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0390= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0390= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0390= (i + 390) % 2;  // Phase3: 翻转
          end
        end

        // pi0391: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0391= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0391= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0391= (i + 391) % 2;  // Phase3: 翻转
          end
        end

        // pi0392: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0392= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0392= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0392= (i + 392) % 2;  // Phase3: 翻转
          end
        end

        // pi0393: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0393= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0393= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0393= (i + 393) % 2;  // Phase3: 翻转
          end
        end

        // pi0394: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0394= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0394= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0394= (i + 394) % 2;  // Phase3: 翻转
          end
        end

        // pi0395: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0395= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0395= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0395= (i + 395) % 2;  // Phase3: 翻转
          end
        end

        // pi0396: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0396= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0396= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0396= (i + 396) % 2;  // Phase3: 翻转
          end
        end

        // pi0397: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0397= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0397= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0397= (i + 397) % 2;  // Phase3: 翻转
          end
        end

        // pi0398: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0398= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0398= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0398= (i + 398) % 2;  // Phase3: 翻转
          end
        end

        // pi0399: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0399= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0399= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0399= (i + 399) % 2;  // Phase3: 翻转
          end
        end

        // pi0400: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0400= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0400= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0400= (i + 400) % 2;  // Phase3: 翻转
          end
        end

        // pi0401: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0401= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0401= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0401= (i + 401) % 2;  // Phase3: 翻转
          end
        end

        // pi0402: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0402= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0402= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0402= (i + 402) % 2;  // Phase3: 翻转
          end
        end

        // pi0403: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0403= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0403= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0403= (i + 403) % 2;  // Phase3: 翻转
          end
        end

        // pi0404: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0404= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0404= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0404= (i + 404) % 2;  // Phase3: 翻转
          end
        end

        // pi0405: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0405= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0405= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0405= (i + 405) % 2;  // Phase3: 翻转
          end
        end

        // pi0406: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0406= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0406= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0406= (i + 406) % 2;  // Phase3: 翻转
          end
        end

        // pi0407: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0407= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0407= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0407= (i + 407) % 2;  // Phase3: 翻转
          end
        end

        // pi0408: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0408= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0408= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0408= (i + 408) % 2;  // Phase3: 翻转
          end
        end

        // pi0409: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0409= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0409= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0409= (i + 409) % 2;  // Phase3: 翻转
          end
        end

        // pi0410: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0410= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0410= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0410= (i + 410) % 2;  // Phase3: 翻转
          end
        end

        // pi0411: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0411= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0411= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0411= (i + 411) % 2;  // Phase3: 翻转
          end
        end

        // pi0412: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0412= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0412= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0412= (i + 412) % 2;  // Phase3: 翻转
          end
        end

        // pi0413: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0413= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0413= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0413= (i + 413) % 2;  // Phase3: 翻转
          end
        end

        // pi0414: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0414= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0414= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0414= (i + 414) % 2;  // Phase3: 翻转
          end
        end

        // pi0415: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0415= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0415= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0415= (i + 415) % 2;  // Phase3: 翻转
          end
        end

        // pi0416: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0416= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0416= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0416= (i + 416) % 2;  // Phase3: 翻转
          end
        end

        // pi0417: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0417= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0417= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0417= (i + 417) % 2;  // Phase3: 翻转
          end
        end

        // pi0418: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0418= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0418= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0418= (i + 418) % 2;  // Phase3: 翻转
          end
        end

        // pi0419: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0419= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0419= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0419= (i + 419) % 2;  // Phase3: 翻转
          end
        end

        // pi0420: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0420= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0420= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0420= (i + 420) % 2;  // Phase3: 翻转
          end
        end

        // pi0421: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0421= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0421= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0421= (i + 421) % 2;  // Phase3: 翻转
          end
        end

        // pi0422: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0422= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0422= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0422= (i + 422) % 2;  // Phase3: 翻转
          end
        end

        // pi0423: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0423= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0423= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0423= (i + 423) % 2;  // Phase3: 翻转
          end
        end

        // pi0424: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0424= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0424= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0424= (i + 424) % 2;  // Phase3: 翻转
          end
        end

        // pi0425: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0425= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0425= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0425= (i + 425) % 2;  // Phase3: 翻转
          end
        end

        // pi0426: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0426= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0426= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0426= (i + 426) % 2;  // Phase3: 翻转
          end
        end

        // pi0427: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0427= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0427= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0427= (i + 427) % 2;  // Phase3: 翻转
          end
        end

        // pi0428: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0428= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0428= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0428= (i + 428) % 2;  // Phase3: 翻转
          end
        end

        // pi0429: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0429= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0429= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0429= (i + 429) % 2;  // Phase3: 翻转
          end
        end

        // pi0430: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0430= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0430= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0430= (i + 430) % 2;  // Phase3: 翻转
          end
        end

        // pi0431: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0431= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0431= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0431= (i + 431) % 2;  // Phase3: 翻转
          end
        end

        // pi0432: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0432= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0432= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0432= (i + 432) % 2;  // Phase3: 翻转
          end
        end

        // pi0433: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0433= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0433= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0433= (i + 433) % 2;  // Phase3: 翻转
          end
        end

        // pi0434: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0434= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0434= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0434= (i + 434) % 2;  // Phase3: 翻转
          end
        end

        // pi0435: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0435= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0435= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0435= (i + 435) % 2;  // Phase3: 翻转
          end
        end

        // pi0436: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0436= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0436= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0436= (i + 436) % 2;  // Phase3: 翻转
          end
        end

        // pi0437: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0437= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0437= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0437= (i + 437) % 2;  // Phase3: 翻转
          end
        end

        // pi0438: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0438= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0438= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0438= (i + 438) % 2;  // Phase3: 翻转
          end
        end

        // pi0439: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0439= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0439= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0439= (i + 439) % 2;  // Phase3: 翻转
          end
        end

        // pi0440: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0440= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0440= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0440= (i + 440) % 2;  // Phase3: 翻转
          end
        end

        // pi0441: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0441= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0441= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0441= (i + 441) % 2;  // Phase3: 翻转
          end
        end

        // pi0442: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0442= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0442= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0442= (i + 442) % 2;  // Phase3: 翻转
          end
        end

        // pi0443: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0443= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0443= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0443= (i + 443) % 2;  // Phase3: 翻转
          end
        end

        // pi0444: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0444= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0444= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0444= (i + 444) % 2;  // Phase3: 翻转
          end
        end

        // pi0445: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0445= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0445= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0445= (i + 445) % 2;  // Phase3: 翻转
          end
        end

        // pi0446: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0446= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0446= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0446= (i + 446) % 2;  // Phase3: 翻转
          end
        end

        // pi0447: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0447= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0447= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0447= (i + 447) % 2;  // Phase3: 翻转
          end
        end

        // pi0448: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0448= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0448= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0448= (i + 448) % 2;  // Phase3: 翻转
          end
        end

        // pi0449: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0449= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0449= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0449= (i + 449) % 2;  // Phase3: 翻转
          end
        end

        // pi0450: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0450= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0450= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0450= (i + 450) % 2;  // Phase3: 翻转
          end
        end

        // pi0451: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0451= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0451= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0451= (i + 451) % 2;  // Phase3: 翻转
          end
        end

        // pi0452: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0452= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0452= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0452= (i + 452) % 2;  // Phase3: 翻转
          end
        end

        // pi0453: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0453= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0453= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0453= (i + 453) % 2;  // Phase3: 翻转
          end
        end

        // pi0454: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0454= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0454= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0454= (i + 454) % 2;  // Phase3: 翻转
          end
        end

        // pi0455: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0455= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0455= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0455= (i + 455) % 2;  // Phase3: 翻转
          end
        end

        // pi0456: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0456= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0456= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0456= (i + 456) % 2;  // Phase3: 翻转
          end
        end

        // pi0457: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0457= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0457= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0457= (i + 457) % 2;  // Phase3: 翻转
          end
        end

        // pi0458: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0458= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0458= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0458= (i + 458) % 2;  // Phase3: 翻转
          end
        end

        // pi0459: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0459= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0459= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0459= (i + 459) % 2;  // Phase3: 翻转
          end
        end

        // pi0460: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0460= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0460= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0460= (i + 460) % 2;  // Phase3: 翻转
          end
        end

        // pi0461: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0461= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0461= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0461= (i + 461) % 2;  // Phase3: 翻转
          end
        end

        // pi0462: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0462= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0462= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0462= (i + 462) % 2;  // Phase3: 翻转
          end
        end

        // pi0463: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0463= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0463= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0463= (i + 463) % 2;  // Phase3: 翻转
          end
        end

        // pi0464: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0464= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0464= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0464= (i + 464) % 2;  // Phase3: 翻转
          end
        end

        // pi0465: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0465= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0465= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0465= (i + 465) % 2;  // Phase3: 翻转
          end
        end

        // pi0466: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0466= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0466= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0466= (i + 466) % 2;  // Phase3: 翻转
          end
        end

        // pi0467: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0467= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0467= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0467= (i + 467) % 2;  // Phase3: 翻转
          end
        end

        // pi0468: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0468= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0468= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0468= (i + 468) % 2;  // Phase3: 翻转
          end
        end

        // pi0469: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0469= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0469= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0469= (i + 469) % 2;  // Phase3: 翻转
          end
        end

        // pi0470: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0470= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0470= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0470= (i + 470) % 2;  // Phase3: 翻转
          end
        end

        // pi0471: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0471= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0471= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0471= (i + 471) % 2;  // Phase3: 翻转
          end
        end

        // pi0472: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0472= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0472= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0472= (i + 472) % 2;  // Phase3: 翻转
          end
        end

        // pi0473: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0473= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0473= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0473= (i + 473) % 2;  // Phase3: 翻转
          end
        end

        // pi0474: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0474= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0474= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0474= (i + 474) % 2;  // Phase3: 翻转
          end
        end

        // pi0475: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0475= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0475= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0475= (i + 475) % 2;  // Phase3: 翻转
          end
        end

        // pi0476: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0476= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0476= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0476= (i + 476) % 2;  // Phase3: 翻转
          end
        end

        // pi0477: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0477= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0477= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0477= (i + 477) % 2;  // Phase3: 翻转
          end
        end

        // pi0478: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0478= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0478= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0478= (i + 478) % 2;  // Phase3: 翻转
          end
        end

        // pi0479: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0479= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0479= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0479= (i + 479) % 2;  // Phase3: 翻转
          end
        end

        // pi0480: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0480= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0480= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0480= (i + 480) % 2;  // Phase3: 翻转
          end
        end

        // pi0481: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0481= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0481= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0481= (i + 481) % 2;  // Phase3: 翻转
          end
        end

        // pi0482: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0482= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0482= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0482= (i + 482) % 2;  // Phase3: 翻转
          end
        end

        // pi0483: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0483= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0483= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0483= (i + 483) % 2;  // Phase3: 翻转
          end
        end

        // pi0484: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0484= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0484= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0484= (i + 484) % 2;  // Phase3: 翻转
          end
        end

        // pi0485: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0485= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0485= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0485= (i + 485) % 2;  // Phase3: 翻转
          end
        end

        // pi0486: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0486= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0486= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0486= (i + 486) % 2;  // Phase3: 翻转
          end
        end

        // pi0487: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0487= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0487= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0487= (i + 487) % 2;  // Phase3: 翻转
          end
        end

        // pi0488: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0488= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0488= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0488= (i + 488) % 2;  // Phase3: 翻转
          end
        end

        // pi0489: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0489= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0489= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0489= (i + 489) % 2;  // Phase3: 翻转
          end
        end

        // pi0490: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0490= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0490= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0490= (i + 490) % 2;  // Phase3: 翻转
          end
        end

        // pi0491: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0491= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0491= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0491= (i + 491) % 2;  // Phase3: 翻转
          end
        end

        // pi0492: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0492= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0492= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0492= (i + 492) % 2;  // Phase3: 翻转
          end
        end

        // pi0493: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0493= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0493= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0493= (i + 493) % 2;  // Phase3: 翻转
          end
        end

        // pi0494: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0494= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0494= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0494= (i + 494) % 2;  // Phase3: 翻转
          end
        end

        // pi0495: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0495= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0495= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0495= (i + 495) % 2;  // Phase3: 翻转
          end
        end

        // pi0496: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0496= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0496= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0496= (i + 496) % 2;  // Phase3: 翻转
          end
        end

        // pi0497: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0497= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0497= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0497= (i + 497) % 2;  // Phase3: 翻转
          end
        end

        // pi0498: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0498= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0498= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0498= (i + 498) % 2;  // Phase3: 翻转
          end
        end

        // pi0499: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0499= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0499= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0499= (i + 499) % 2;  // Phase3: 翻转
          end
        end

        // pi0500: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0500= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0500= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0500= (i + 500) % 2;  // Phase3: 翻转
          end
        end

        // pi0501: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0501= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0501= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0501= (i + 501) % 2;  // Phase3: 翻转
          end
        end

        // pi0502: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0502= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0502= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0502= (i + 502) % 2;  // Phase3: 翻转
          end
        end

        // pi0503: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0503= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0503= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0503= (i + 503) % 2;  // Phase3: 翻转
          end
        end

        // pi0504: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0504= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0504= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0504= (i + 504) % 2;  // Phase3: 翻转
          end
        end

        // pi0505: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0505= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0505= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0505= (i + 505) % 2;  // Phase3: 翻转
          end
        end

        // pi0506: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0506= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0506= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0506= (i + 506) % 2;  // Phase3: 翻转
          end
        end

        // pi0507: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0507= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0507= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0507= (i + 507) % 2;  // Phase3: 翻转
          end
        end

        // pi0508: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0508= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0508= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0508= (i + 508) % 2;  // Phase3: 翻转
          end
        end

        // pi0509: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0509= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0509= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0509= (i + 509) % 2;  // Phase3: 翻转
          end
        end

        // pi0510: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0510= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0510= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0510= (i + 510) % 2;  // Phase3: 翻转
          end
        end

        // pi0511: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0511= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0511= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0511= (i + 511) % 2;  // Phase3: 翻转
          end
        end

        // pi0512: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0512= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0512= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0512= (i + 512) % 2;  // Phase3: 翻转
          end
        end

        // pi0513: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0513= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0513= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0513= (i + 513) % 2;  // Phase3: 翻转
          end
        end

        // pi0514: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0514= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0514= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0514= (i + 514) % 2;  // Phase3: 翻转
          end
        end

        // pi0515: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0515= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0515= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0515= (i + 515) % 2;  // Phase3: 翻转
          end
        end

        // pi0516: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0516= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0516= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0516= (i + 516) % 2;  // Phase3: 翻转
          end
        end

        // pi0517: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0517= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0517= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0517= (i + 517) % 2;  // Phase3: 翻转
          end
        end

        // pi0518: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0518= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0518= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0518= (i + 518) % 2;  // Phase3: 翻转
          end
        end

        // pi0519: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0519= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0519= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0519= (i + 519) % 2;  // Phase3: 翻转
          end
        end

        // pi0520: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0520= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0520= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0520= (i + 520) % 2;  // Phase3: 翻转
          end
        end

        // pi0521: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0521= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0521= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0521= (i + 521) % 2;  // Phase3: 翻转
          end
        end

        // pi0522: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0522= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0522= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0522= (i + 522) % 2;  // Phase3: 翻转
          end
        end

        // pi0523: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0523= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0523= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0523= (i + 523) % 2;  // Phase3: 翻转
          end
        end

        // pi0524: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0524= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0524= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0524= (i + 524) % 2;  // Phase3: 翻转
          end
        end

        // pi0525: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0525= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0525= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0525= (i + 525) % 2;  // Phase3: 翻转
          end
        end

        // pi0526: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0526= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0526= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0526= (i + 526) % 2;  // Phase3: 翻转
          end
        end

        // pi0527: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0527= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0527= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0527= (i + 527) % 2;  // Phase3: 翻转
          end
        end

        // pi0528: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0528= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0528= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0528= (i + 528) % 2;  // Phase3: 翻转
          end
        end

        // pi0529: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0529= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0529= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0529= (i + 529) % 2;  // Phase3: 翻转
          end
        end

        // pi0530: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0530= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0530= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0530= (i + 530) % 2;  // Phase3: 翻转
          end
        end

        // pi0531: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0531= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0531= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0531= (i + 531) % 2;  // Phase3: 翻转
          end
        end

        // pi0532: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0532= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0532= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0532= (i + 532) % 2;  // Phase3: 翻转
          end
        end

        // pi0533: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0533= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0533= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0533= (i + 533) % 2;  // Phase3: 翻转
          end
        end

        // pi0534: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0534= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0534= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0534= (i + 534) % 2;  // Phase3: 翻转
          end
        end

        // pi0535: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0535= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0535= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0535= (i + 535) % 2;  // Phase3: 翻转
          end
        end

        // pi0536: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0536= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0536= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0536= (i + 536) % 2;  // Phase3: 翻转
          end
        end

        // pi0537: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0537= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0537= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0537= (i + 537) % 2;  // Phase3: 翻转
          end
        end

        // pi0538: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0538= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0538= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0538= (i + 538) % 2;  // Phase3: 翻转
          end
        end

        // pi0539: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0539= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0539= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0539= (i + 539) % 2;  // Phase3: 翻转
          end
        end

        // pi0540: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0540= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0540= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0540= (i + 540) % 2;  // Phase3: 翻转
          end
        end

        // pi0541: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0541= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0541= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0541= (i + 541) % 2;  // Phase3: 翻转
          end
        end

        // pi0542: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0542= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0542= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0542= (i + 542) % 2;  // Phase3: 翻转
          end
        end

        // pi0543: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0543= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0543= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0543= (i + 543) % 2;  // Phase3: 翻转
          end
        end

        // pi0544: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0544= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0544= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0544= (i + 544) % 2;  // Phase3: 翻转
          end
        end

        // pi0545: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0545= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0545= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0545= (i + 545) % 2;  // Phase3: 翻转
          end
        end

        // pi0546: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0546= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0546= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0546= (i + 546) % 2;  // Phase3: 翻转
          end
        end

        // pi0547: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0547= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0547= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0547= (i + 547) % 2;  // Phase3: 翻转
          end
        end

        // pi0548: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0548= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0548= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0548= (i + 548) % 2;  // Phase3: 翻转
          end
        end

        // pi0549: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0549= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0549= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0549= (i + 549) % 2;  // Phase3: 翻转
          end
        end

        // pi0550: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0550= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0550= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0550= (i + 550) % 2;  // Phase3: 翻转
          end
        end

        // pi0551: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0551= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0551= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0551= (i + 551) % 2;  // Phase3: 翻转
          end
        end

        // pi0552: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0552= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0552= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0552= (i + 552) % 2;  // Phase3: 翻转
          end
        end

        // pi0553: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0553= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0553= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0553= (i + 553) % 2;  // Phase3: 翻转
          end
        end

        // pi0554: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0554= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0554= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0554= (i + 554) % 2;  // Phase3: 翻转
          end
        end

        // pi0555: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0555= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0555= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0555= (i + 555) % 2;  // Phase3: 翻转
          end
        end

        // pi0556: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0556= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0556= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0556= (i + 556) % 2;  // Phase3: 翻转
          end
        end

        // pi0557: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0557= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0557= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0557= (i + 557) % 2;  // Phase3: 翻转
          end
        end

        // pi0558: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0558= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0558= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0558= (i + 558) % 2;  // Phase3: 翻转
          end
        end

        // pi0559: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0559= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0559= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0559= (i + 559) % 2;  // Phase3: 翻转
          end
        end

        // pi0560: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0560= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0560= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0560= (i + 560) % 2;  // Phase3: 翻转
          end
        end

        // pi0561: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0561= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0561= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0561= (i + 561) % 2;  // Phase3: 翻转
          end
        end

        // pi0562: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0562= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0562= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0562= (i + 562) % 2;  // Phase3: 翻转
          end
        end

        // pi0563: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0563= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0563= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0563= (i + 563) % 2;  // Phase3: 翻转
          end
        end

        // pi0564: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0564= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0564= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0564= (i + 564) % 2;  // Phase3: 翻转
          end
        end

        // pi0565: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0565= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0565= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0565= (i + 565) % 2;  // Phase3: 翻转
          end
        end

        // pi0566: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0566= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0566= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0566= (i + 566) % 2;  // Phase3: 翻转
          end
        end

        // pi0567: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0567= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0567= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0567= (i + 567) % 2;  // Phase3: 翻转
          end
        end

        // pi0568: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0568= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0568= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0568= (i + 568) % 2;  // Phase3: 翻转
          end
        end

        // pi0569: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0569= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0569= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0569= (i + 569) % 2;  // Phase3: 翻转
          end
        end

        // pi0570: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0570= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0570= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0570= (i + 570) % 2;  // Phase3: 翻转
          end
        end

        // pi0571: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0571= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0571= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0571= (i + 571) % 2;  // Phase3: 翻转
          end
        end

        // pi0572: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0572= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0572= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0572= (i + 572) % 2;  // Phase3: 翻转
          end
        end

        // pi0573: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0573= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0573= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0573= (i + 573) % 2;  // Phase3: 翻转
          end
        end

        // pi0574: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0574= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0574= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0574= (i + 574) % 2;  // Phase3: 翻转
          end
        end

        // pi0575: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0575= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0575= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0575= (i + 575) % 2;  // Phase3: 翻转
          end
        end

        // pi0576: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0576= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0576= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0576= (i + 576) % 2;  // Phase3: 翻转
          end
        end

        // pi0577: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0577= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0577= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0577= (i + 577) % 2;  // Phase3: 翻转
          end
        end

        // pi0578: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0578= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0578= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0578= (i + 578) % 2;  // Phase3: 翻转
          end
        end

        // pi0579: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0579= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0579= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0579= (i + 579) % 2;  // Phase3: 翻转
          end
        end

        // pi0580: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0580= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0580= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0580= (i + 580) % 2;  // Phase3: 翻转
          end
        end

        // pi0581: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0581= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0581= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0581= (i + 581) % 2;  // Phase3: 翻转
          end
        end

        // pi0582: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0582= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0582= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0582= (i + 582) % 2;  // Phase3: 翻转
          end
        end

        // pi0583: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0583= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0583= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0583= (i + 583) % 2;  // Phase3: 翻转
          end
        end

        // pi0584: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0584= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0584= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0584= (i + 584) % 2;  // Phase3: 翻转
          end
        end

        // pi0585: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0585= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0585= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0585= (i + 585) % 2;  // Phase3: 翻转
          end
        end

        // pi0586: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0586= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0586= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0586= (i + 586) % 2;  // Phase3: 翻转
          end
        end

        // pi0587: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0587= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0587= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0587= (i + 587) % 2;  // Phase3: 翻转
          end
        end

        // pi0588: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0588= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0588= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0588= (i + 588) % 2;  // Phase3: 翻转
          end
        end

        // pi0589: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0589= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0589= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0589= (i + 589) % 2;  // Phase3: 翻转
          end
        end

        // pi0590: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0590= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0590= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0590= (i + 590) % 2;  // Phase3: 翻转
          end
        end

        // pi0591: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0591= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0591= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0591= (i + 591) % 2;  // Phase3: 翻转
          end
        end

        // pi0592: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0592= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0592= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0592= (i + 592) % 2;  // Phase3: 翻转
          end
        end

        // pi0593: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0593= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0593= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0593= (i + 593) % 2;  // Phase3: 翻转
          end
        end

        // pi0594: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0594= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0594= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0594= (i + 594) % 2;  // Phase3: 翻转
          end
        end

        // pi0595: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0595= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0595= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0595= (i + 595) % 2;  // Phase3: 翻转
          end
        end

        // pi0596: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0596= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0596= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0596= (i + 596) % 2;  // Phase3: 翻转
          end
        end

        // pi0597: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0597= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0597= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0597= (i + 597) % 2;  // Phase3: 翻转
          end
        end

        // pi0598: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0598= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0598= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0598= (i + 598) % 2;  // Phase3: 翻转
          end
        end

        // pi0599: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0599= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0599= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0599= (i + 599) % 2;  // Phase3: 翻转
          end
        end

        // pi0600: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0600= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0600= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0600= (i + 600) % 2;  // Phase3: 翻转
          end
        end

        // pi0601: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0601= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0601= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0601= (i + 601) % 2;  // Phase3: 翻转
          end
        end

        // pi0602: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0602= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0602= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0602= (i + 602) % 2;  // Phase3: 翻转
          end
        end

        // pi0603: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0603= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0603= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0603= (i + 603) % 2;  // Phase3: 翻转
          end
        end

        // pi0604: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0604= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0604= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0604= (i + 604) % 2;  // Phase3: 翻转
          end
        end

        // pi0605: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0605= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0605= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0605= (i + 605) % 2;  // Phase3: 翻转
          end
        end

        // pi0606: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0606= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0606= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0606= (i + 606) % 2;  // Phase3: 翻转
          end
        end

        // pi0607: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0607= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0607= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0607= (i + 607) % 2;  // Phase3: 翻转
          end
        end

        // pi0608: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0608= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0608= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0608= (i + 608) % 2;  // Phase3: 翻转
          end
        end

        // pi0609: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0609= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0609= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0609= (i + 609) % 2;  // Phase3: 翻转
          end
        end

        // pi0610: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0610= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0610= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0610= (i + 610) % 2;  // Phase3: 翻转
          end
        end

        // pi0611: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0611= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0611= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0611= (i + 611) % 2;  // Phase3: 翻转
          end
        end

        // pi0612: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0612= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0612= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0612= (i + 612) % 2;  // Phase3: 翻转
          end
        end

        // pi0613: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0613= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0613= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0613= (i + 613) % 2;  // Phase3: 翻转
          end
        end

        // pi0614: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0614= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0614= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0614= (i + 614) % 2;  // Phase3: 翻转
          end
        end

        // pi0615: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0615= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0615= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0615= (i + 615) % 2;  // Phase3: 翻转
          end
        end

        // pi0616: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0616= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0616= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0616= (i + 616) % 2;  // Phase3: 翻转
          end
        end

        // pi0617: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0617= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0617= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0617= (i + 617) % 2;  // Phase3: 翻转
          end
        end

        // pi0618: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0618= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0618= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0618= (i + 618) % 2;  // Phase3: 翻转
          end
        end

        // pi0619: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0619= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0619= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0619= (i + 619) % 2;  // Phase3: 翻转
          end
        end

        // pi0620: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0620= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0620= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0620= (i + 620) % 2;  // Phase3: 翻转
          end
        end

        // pi0621: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0621= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0621= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0621= (i + 621) % 2;  // Phase3: 翻转
          end
        end

        // pi0622: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0622= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0622= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0622= (i + 622) % 2;  // Phase3: 翻转
          end
        end

        // pi0623: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0623= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0623= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0623= (i + 623) % 2;  // Phase3: 翻转
          end
        end

        // pi0624: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0624= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0624= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0624= (i + 624) % 2;  // Phase3: 翻转
          end
        end

        // pi0625: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0625= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0625= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0625= (i + 625) % 2;  // Phase3: 翻转
          end
        end

        // pi0626: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0626= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0626= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0626= (i + 626) % 2;  // Phase3: 翻转
          end
        end

        // pi0627: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0627= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0627= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0627= (i + 627) % 2;  // Phase3: 翻转
          end
        end

        // pi0628: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0628= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0628= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0628= (i + 628) % 2;  // Phase3: 翻转
          end
        end

        // pi0629: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0629= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0629= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0629= (i + 629) % 2;  // Phase3: 翻转
          end
        end

        // pi0630: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0630= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0630= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0630= (i + 630) % 2;  // Phase3: 翻转
          end
        end

        // pi0631: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0631= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0631= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0631= (i + 631) % 2;  // Phase3: 翻转
          end
        end

        // pi0632: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0632= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0632= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0632= (i + 632) % 2;  // Phase3: 翻转
          end
        end

        // pi0633: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0633= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0633= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0633= (i + 633) % 2;  // Phase3: 翻转
          end
        end

        // pi0634: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0634= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0634= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0634= (i + 634) % 2;  // Phase3: 翻转
          end
        end

        // pi0635: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0635= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0635= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0635= (i + 635) % 2;  // Phase3: 翻转
          end
        end

        // pi0636: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0636= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0636= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0636= (i + 636) % 2;  // Phase3: 翻转
          end
        end

        // pi0637: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0637= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0637= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0637= (i + 637) % 2;  // Phase3: 翻转
          end
        end

        // pi0638: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0638= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0638= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0638= (i + 638) % 2;  // Phase3: 翻转
          end
        end

        // pi0639: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0639= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0639= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0639= (i + 639) % 2;  // Phase3: 翻转
          end
        end

        // pi0640: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0640= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0640= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0640= (i + 640) % 2;  // Phase3: 翻转
          end
        end

        // pi0641: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0641= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0641= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0641= (i + 641) % 2;  // Phase3: 翻转
          end
        end

        // pi0642: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0642= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0642= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0642= (i + 642) % 2;  // Phase3: 翻转
          end
        end

        // pi0643: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0643= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0643= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0643= (i + 643) % 2;  // Phase3: 翻转
          end
        end

        // pi0644: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0644= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0644= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0644= (i + 644) % 2;  // Phase3: 翻转
          end
        end

        // pi0645: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0645= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0645= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0645= (i + 645) % 2;  // Phase3: 翻转
          end
        end

        // pi0646: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0646= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0646= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0646= (i + 646) % 2;  // Phase3: 翻转
          end
        end

        // pi0647: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0647= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0647= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0647= (i + 647) % 2;  // Phase3: 翻转
          end
        end

        // pi0648: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0648= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0648= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0648= (i + 648) % 2;  // Phase3: 翻转
          end
        end

        // pi0649: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0649= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0649= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0649= (i + 649) % 2;  // Phase3: 翻转
          end
        end

        // pi0650: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0650= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0650= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0650= (i + 650) % 2;  // Phase3: 翻转
          end
        end

        // pi0651: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0651= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0651= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0651= (i + 651) % 2;  // Phase3: 翻转
          end
        end

        // pi0652: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0652= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0652= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0652= (i + 652) % 2;  // Phase3: 翻转
          end
        end

        // pi0653: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0653= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0653= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0653= (i + 653) % 2;  // Phase3: 翻转
          end
        end

        // pi0654: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0654= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0654= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0654= (i + 654) % 2;  // Phase3: 翻转
          end
        end

        // pi0655: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0655= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0655= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0655= (i + 655) % 2;  // Phase3: 翻转
          end
        end

        // pi0656: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0656= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0656= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0656= (i + 656) % 2;  // Phase3: 翻转
          end
        end

        // pi0657: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0657= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0657= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0657= (i + 657) % 2;  // Phase3: 翻转
          end
        end

        // pi0658: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0658= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0658= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0658= (i + 658) % 2;  // Phase3: 翻转
          end
        end

        // pi0659: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0659= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0659= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0659= (i + 659) % 2;  // Phase3: 翻转
          end
        end

        // pi0660: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0660= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0660= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0660= (i + 660) % 2;  // Phase3: 翻转
          end
        end

        // pi0661: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0661= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0661= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0661= (i + 661) % 2;  // Phase3: 翻转
          end
        end

        // pi0662: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0662= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0662= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0662= (i + 662) % 2;  // Phase3: 翻转
          end
        end

        // pi0663: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0663= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0663= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0663= (i + 663) % 2;  // Phase3: 翻转
          end
        end

        // pi0664: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0664= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0664= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0664= (i + 664) % 2;  // Phase3: 翻转
          end
        end

        // pi0665: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0665= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0665= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0665= (i + 665) % 2;  // Phase3: 翻转
          end
        end

        // pi0666: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0666= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0666= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0666= (i + 666) % 2;  // Phase3: 翻转
          end
        end

        // pi0667: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0667= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0667= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0667= (i + 667) % 2;  // Phase3: 翻转
          end
        end

        // pi0668: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0668= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0668= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0668= (i + 668) % 2;  // Phase3: 翻转
          end
        end

        // pi0669: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0669= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0669= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0669= (i + 669) % 2;  // Phase3: 翻转
          end
        end

        // pi0670: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0670= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0670= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0670= (i + 670) % 2;  // Phase3: 翻转
          end
        end

        // pi0671: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0671= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0671= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0671= (i + 671) % 2;  // Phase3: 翻转
          end
        end

        // pi0672: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0672= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0672= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0672= (i + 672) % 2;  // Phase3: 翻转
          end
        end

        // pi0673: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0673= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0673= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0673= (i + 673) % 2;  // Phase3: 翻转
          end
        end

        // pi0674: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0674= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0674= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0674= (i + 674) % 2;  // Phase3: 翻转
          end
        end

        // pi0675: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0675= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0675= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0675= (i + 675) % 2;  // Phase3: 翻转
          end
        end

        // pi0676: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0676= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0676= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0676= (i + 676) % 2;  // Phase3: 翻转
          end
        end

        // pi0677: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0677= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0677= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0677= (i + 677) % 2;  // Phase3: 翻转
          end
        end

        // pi0678: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0678= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0678= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0678= (i + 678) % 2;  // Phase3: 翻转
          end
        end

        // pi0679: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0679= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0679= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0679= (i + 679) % 2;  // Phase3: 翻转
          end
        end

        // pi0680: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0680= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0680= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0680= (i + 680) % 2;  // Phase3: 翻转
          end
        end

        // pi0681: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0681= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0681= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0681= (i + 681) % 2;  // Phase3: 翻转
          end
        end

        // pi0682: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0682= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0682= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0682= (i + 682) % 2;  // Phase3: 翻转
          end
        end

        // pi0683: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0683= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0683= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0683= (i + 683) % 2;  // Phase3: 翻转
          end
        end

        // pi0684: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0684= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0684= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0684= (i + 684) % 2;  // Phase3: 翻转
          end
        end

        // pi0685: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0685= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0685= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0685= (i + 685) % 2;  // Phase3: 翻转
          end
        end

        // pi0686: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0686= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0686= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0686= (i + 686) % 2;  // Phase3: 翻转
          end
        end

        // pi0687: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0687= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0687= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0687= (i + 687) % 2;  // Phase3: 翻转
          end
        end

        // pi0688: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0688= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0688= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0688= (i + 688) % 2;  // Phase3: 翻转
          end
        end

        // pi0689: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0689= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0689= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0689= (i + 689) % 2;  // Phase3: 翻转
          end
        end

        // pi0690: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0690= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0690= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0690= (i + 690) % 2;  // Phase3: 翻转
          end
        end

        // pi0691: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0691= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0691= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0691= (i + 691) % 2;  // Phase3: 翻转
          end
        end

        // pi0692: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0692= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0692= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0692= (i + 692) % 2;  // Phase3: 翻转
          end
        end

        // pi0693: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0693= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0693= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0693= (i + 693) % 2;  // Phase3: 翻转
          end
        end

        // pi0694: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0694= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0694= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0694= (i + 694) % 2;  // Phase3: 翻转
          end
        end

        // pi0695: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0695= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0695= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0695= (i + 695) % 2;  // Phase3: 翻转
          end
        end

        // pi0696: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0696= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0696= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0696= (i + 696) % 2;  // Phase3: 翻转
          end
        end

        // pi0697: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0697= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0697= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0697= (i + 697) % 2;  // Phase3: 翻转
          end
        end

        // pi0698: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0698= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0698= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0698= (i + 698) % 2;  // Phase3: 翻转
          end
        end

        // pi0699: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0699= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0699= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0699= (i + 699) % 2;  // Phase3: 翻转
          end
        end

        // pi0700: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0700= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0700= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0700= (i + 700) % 2;  // Phase3: 翻转
          end
        end

        // pi0701: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0701= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0701= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0701= (i + 701) % 2;  // Phase3: 翻转
          end
        end

        // pi0702: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0702= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0702= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0702= (i + 702) % 2;  // Phase3: 翻转
          end
        end

        // pi0703: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0703= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0703= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0703= (i + 703) % 2;  // Phase3: 翻转
          end
        end

        // pi0704: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0704= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0704= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0704= (i + 704) % 2;  // Phase3: 翻转
          end
        end

        // pi0705: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0705= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0705= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0705= (i + 705) % 2;  // Phase3: 翻转
          end
        end

        // pi0706: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0706= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0706= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0706= (i + 706) % 2;  // Phase3: 翻转
          end
        end

        // pi0707: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0707= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0707= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0707= (i + 707) % 2;  // Phase3: 翻转
          end
        end

        // pi0708: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0708= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0708= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0708= (i + 708) % 2;  // Phase3: 翻转
          end
        end

        // pi0709: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0709= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0709= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0709= (i + 709) % 2;  // Phase3: 翻转
          end
        end

        // pi0710: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0710= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0710= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0710= (i + 710) % 2;  // Phase3: 翻转
          end
        end

        // pi0711: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0711= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0711= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0711= (i + 711) % 2;  // Phase3: 翻转
          end
        end

        // pi0712: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0712= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0712= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0712= (i + 712) % 2;  // Phase3: 翻转
          end
        end

        // pi0713: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0713= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0713= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0713= (i + 713) % 2;  // Phase3: 翻转
          end
        end

        // pi0714: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0714= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0714= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0714= (i + 714) % 2;  // Phase3: 翻转
          end
        end

        // pi0715: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0715= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0715= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0715= (i + 715) % 2;  // Phase3: 翻转
          end
        end

        // pi0716: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0716= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0716= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0716= (i + 716) % 2;  // Phase3: 翻转
          end
        end

        // pi0717: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0717= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0717= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0717= (i + 717) % 2;  // Phase3: 翻转
          end
        end

        // pi0718: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0718= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0718= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0718= (i + 718) % 2;  // Phase3: 翻转
          end
        end

        // pi0719: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0719= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0719= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0719= (i + 719) % 2;  // Phase3: 翻转
          end
        end

        // pi0720: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0720= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0720= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0720= (i + 720) % 2;  // Phase3: 翻转
          end
        end

        // pi0721: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0721= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0721= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0721= (i + 721) % 2;  // Phase3: 翻转
          end
        end

        // pi0722: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0722= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0722= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0722= (i + 722) % 2;  // Phase3: 翻转
          end
        end

        // pi0723: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0723= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0723= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0723= (i + 723) % 2;  // Phase3: 翻转
          end
        end

        // pi0724: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0724= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0724= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0724= (i + 724) % 2;  // Phase3: 翻转
          end
        end

        // pi0725: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0725= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0725= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0725= (i + 725) % 2;  // Phase3: 翻转
          end
        end

        // pi0726: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0726= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0726= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0726= (i + 726) % 2;  // Phase3: 翻转
          end
        end

        // pi0727: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0727= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0727= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0727= (i + 727) % 2;  // Phase3: 翻转
          end
        end

        // pi0728: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0728= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0728= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0728= (i + 728) % 2;  // Phase3: 翻转
          end
        end

        // pi0729: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0729= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0729= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0729= (i + 729) % 2;  // Phase3: 翻转
          end
        end

        // pi0730: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0730= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0730= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0730= (i + 730) % 2;  // Phase3: 翻转
          end
        end

        // pi0731: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0731= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0731= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0731= (i + 731) % 2;  // Phase3: 翻转
          end
        end

        // pi0732: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0732= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0732= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0732= (i + 732) % 2;  // Phase3: 翻转
          end
        end

        // pi0733: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0733= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0733= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0733= (i + 733) % 2;  // Phase3: 翻转
          end
        end

        // pi0734: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0734= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0734= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0734= (i + 734) % 2;  // Phase3: 翻转
          end
        end

        // pi0735: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0735= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0735= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0735= (i + 735) % 2;  // Phase3: 翻转
          end
        end

        // pi0736: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0736= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0736= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0736= (i + 736) % 2;  // Phase3: 翻转
          end
        end

        // pi0737: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0737= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0737= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0737= (i + 737) % 2;  // Phase3: 翻转
          end
        end

        // pi0738: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0738= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0738= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0738= (i + 738) % 2;  // Phase3: 翻转
          end
        end

        // pi0739: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0739= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0739= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0739= (i + 739) % 2;  // Phase3: 翻转
          end
        end

        // pi0740: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0740= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0740= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0740= (i + 740) % 2;  // Phase3: 翻转
          end
        end

        // pi0741: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0741= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0741= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0741= (i + 741) % 2;  // Phase3: 翻转
          end
        end

        // pi0742: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0742= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0742= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0742= (i + 742) % 2;  // Phase3: 翻转
          end
        end

        // pi0743: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0743= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0743= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0743= (i + 743) % 2;  // Phase3: 翻转
          end
        end

        // pi0744: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0744= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0744= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0744= (i + 744) % 2;  // Phase3: 翻转
          end
        end

        // pi0745: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0745= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0745= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0745= (i + 745) % 2;  // Phase3: 翻转
          end
        end

        // pi0746: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0746= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0746= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0746= (i + 746) % 2;  // Phase3: 翻转
          end
        end

        // pi0747: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0747= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0747= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0747= (i + 747) % 2;  // Phase3: 翻转
          end
        end

        // pi0748: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0748= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0748= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0748= (i + 748) % 2;  // Phase3: 翻转
          end
        end

        // pi0749: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0749= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0749= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0749= (i + 749) % 2;  // Phase3: 翻转
          end
        end

        // pi0750: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0750= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0750= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0750= (i + 750) % 2;  // Phase3: 翻转
          end
        end

        // pi0751: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0751= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0751= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0751= (i + 751) % 2;  // Phase3: 翻转
          end
        end

        // pi0752: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0752= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0752= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0752= (i + 752) % 2;  // Phase3: 翻转
          end
        end

        // pi0753: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0753= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0753= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0753= (i + 753) % 2;  // Phase3: 翻转
          end
        end

        // pi0754: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0754= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0754= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0754= (i + 754) % 2;  // Phase3: 翻转
          end
        end

        // pi0755: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0755= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0755= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0755= (i + 755) % 2;  // Phase3: 翻转
          end
        end

        // pi0756: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0756= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0756= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0756= (i + 756) % 2;  // Phase3: 翻转
          end
        end

        // pi0757: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0757= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0757= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0757= (i + 757) % 2;  // Phase3: 翻转
          end
        end

        // pi0758: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0758= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0758= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0758= (i + 758) % 2;  // Phase3: 翻转
          end
        end

        // pi0759: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0759= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0759= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0759= (i + 759) % 2;  // Phase3: 翻转
          end
        end

        // pi0760: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0760= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0760= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0760= (i + 760) % 2;  // Phase3: 翻转
          end
        end

        // pi0761: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0761= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0761= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0761= (i + 761) % 2;  // Phase3: 翻转
          end
        end

        // pi0762: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0762= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0762= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0762= (i + 762) % 2;  // Phase3: 翻转
          end
        end

        // pi0763: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0763= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0763= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0763= (i + 763) % 2;  // Phase3: 翻转
          end
        end

        // pi0764: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0764= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0764= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0764= (i + 764) % 2;  // Phase3: 翻转
          end
        end

        // pi0765: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0765= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0765= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0765= (i + 765) % 2;  // Phase3: 翻转
          end
        end

        // pi0766: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0766= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0766= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0766= (i + 766) % 2;  // Phase3: 翻转
          end
        end

        // pi0767: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0767= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0767= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0767= (i + 767) % 2;  // Phase3: 翻转
          end
        end

        // pi0768: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0768= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0768= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0768= (i + 768) % 2;  // Phase3: 翻转
          end
        end

        // pi0769: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0769= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0769= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0769= (i + 769) % 2;  // Phase3: 翻转
          end
        end

        // pi0770: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0770= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0770= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0770= (i + 770) % 2;  // Phase3: 翻转
          end
        end

        // pi0771: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0771= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0771= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0771= (i + 771) % 2;  // Phase3: 翻转
          end
        end

        // pi0772: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0772= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0772= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0772= (i + 772) % 2;  // Phase3: 翻转
          end
        end

        // pi0773: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0773= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0773= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0773= (i + 773) % 2;  // Phase3: 翻转
          end
        end

        // pi0774: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0774= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0774= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0774= (i + 774) % 2;  // Phase3: 翻转
          end
        end

        // pi0775: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0775= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0775= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0775= (i + 775) % 2;  // Phase3: 翻转
          end
        end

        // pi0776: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0776= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0776= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0776= (i + 776) % 2;  // Phase3: 翻转
          end
        end

        // pi0777: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0777= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0777= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0777= (i + 777) % 2;  // Phase3: 翻转
          end
        end

        // pi0778: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0778= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0778= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0778= (i + 778) % 2;  // Phase3: 翻转
          end
        end

        // pi0779: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0779= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0779= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0779= (i + 779) % 2;  // Phase3: 翻转
          end
        end

        // pi0780: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0780= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0780= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0780= (i + 780) % 2;  // Phase3: 翻转
          end
        end

        // pi0781: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0781= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0781= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0781= (i + 781) % 2;  // Phase3: 翻转
          end
        end

        // pi0782: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0782= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0782= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0782= (i + 782) % 2;  // Phase3: 翻转
          end
        end

        // pi0783: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0783= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0783= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0783= (i + 783) % 2;  // Phase3: 翻转
          end
        end

        // pi0784: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0784= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0784= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0784= (i + 784) % 2;  // Phase3: 翻转
          end
        end

        // pi0785: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0785= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0785= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0785= (i + 785) % 2;  // Phase3: 翻转
          end
        end

        // pi0786: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0786= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0786= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0786= (i + 786) % 2;  // Phase3: 翻转
          end
        end

        // pi0787: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0787= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0787= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0787= (i + 787) % 2;  // Phase3: 翻转
          end
        end

        // pi0788: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0788= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0788= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0788= (i + 788) % 2;  // Phase3: 翻转
          end
        end

        // pi0789: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0789= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0789= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0789= (i + 789) % 2;  // Phase3: 翻转
          end
        end

        // pi0790: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0790= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0790= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0790= (i + 790) % 2;  // Phase3: 翻转
          end
        end

        // pi0791: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0791= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0791= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0791= (i + 791) % 2;  // Phase3: 翻转
          end
        end

        // pi0792: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0792= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0792= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0792= (i + 792) % 2;  // Phase3: 翻转
          end
        end

        // pi0793: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0793= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0793= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0793= (i + 793) % 2;  // Phase3: 翻转
          end
        end

        // pi0794: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0794= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0794= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0794= (i + 794) % 2;  // Phase3: 翻转
          end
        end

        // pi0795: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0795= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0795= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0795= (i + 795) % 2;  // Phase3: 翻转
          end
        end

        // pi0796: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0796= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0796= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0796= (i + 796) % 2;  // Phase3: 翻转
          end
        end

        // pi0797: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0797= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0797= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0797= (i + 797) % 2;  // Phase3: 翻转
          end
        end

        // pi0798: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0798= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0798= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0798= (i + 798) % 2;  // Phase3: 翻转
          end
        end

        // pi0799: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0799= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0799= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0799= (i + 799) % 2;  // Phase3: 翻转
          end
        end

        // pi0800: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0800= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0800= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0800= (i + 800) % 2;  // Phase3: 翻转
          end
        end

        // pi0801: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0801= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0801= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0801= (i + 801) % 2;  // Phase3: 翻转
          end
        end

        // pi0802: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0802= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0802= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0802= (i + 802) % 2;  // Phase3: 翻转
          end
        end

        // pi0803: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0803= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0803= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0803= (i + 803) % 2;  // Phase3: 翻转
          end
        end

        // pi0804: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0804= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0804= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0804= (i + 804) % 2;  // Phase3: 翻转
          end
        end

        // pi0805: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0805= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0805= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0805= (i + 805) % 2;  // Phase3: 翻转
          end
        end

        // pi0806: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0806= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0806= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0806= (i + 806) % 2;  // Phase3: 翻转
          end
        end

        // pi0807: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0807= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0807= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0807= (i + 807) % 2;  // Phase3: 翻转
          end
        end

        // pi0808: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0808= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0808= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0808= (i + 808) % 2;  // Phase3: 翻转
          end
        end

        // pi0809: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0809= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0809= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0809= (i + 809) % 2;  // Phase3: 翻转
          end
        end

        // pi0810: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0810= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0810= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0810= (i + 810) % 2;  // Phase3: 翻转
          end
        end

        // pi0811: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0811= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0811= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0811= (i + 811) % 2;  // Phase3: 翻转
          end
        end

        // pi0812: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0812= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0812= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0812= (i + 812) % 2;  // Phase3: 翻转
          end
        end

        // pi0813: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0813= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0813= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0813= (i + 813) % 2;  // Phase3: 翻转
          end
        end

        // pi0814: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0814= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0814= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0814= (i + 814) % 2;  // Phase3: 翻转
          end
        end

        // pi0815: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0815= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0815= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0815= (i + 815) % 2;  // Phase3: 翻转
          end
        end

        // pi0816: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0816= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0816= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0816= (i + 816) % 2;  // Phase3: 翻转
          end
        end

        // pi0817: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0817= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0817= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0817= (i + 817) % 2;  // Phase3: 翻转
          end
        end

        // pi0818: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0818= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0818= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0818= (i + 818) % 2;  // Phase3: 翻转
          end
        end

        // pi0819: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0819= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0819= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0819= (i + 819) % 2;  // Phase3: 翻转
          end
        end

        // pi0820: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0820= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0820= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0820= (i + 820) % 2;  // Phase3: 翻转
          end
        end

        // pi0821: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0821= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0821= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0821= (i + 821) % 2;  // Phase3: 翻转
          end
        end

        // pi0822: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0822= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0822= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0822= (i + 822) % 2;  // Phase3: 翻转
          end
        end

        // pi0823: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0823= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0823= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0823= (i + 823) % 2;  // Phase3: 翻转
          end
        end

        // pi0824: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0824= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0824= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0824= (i + 824) % 2;  // Phase3: 翻转
          end
        end

        // pi0825: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0825= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0825= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0825= (i + 825) % 2;  // Phase3: 翻转
          end
        end

        // pi0826: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0826= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0826= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0826= (i + 826) % 2;  // Phase3: 翻转
          end
        end

        // pi0827: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0827= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0827= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0827= (i + 827) % 2;  // Phase3: 翻转
          end
        end

        // pi0828: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0828= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0828= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0828= (i + 828) % 2;  // Phase3: 翻转
          end
        end

        // pi0829: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0829= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0829= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0829= (i + 829) % 2;  // Phase3: 翻转
          end
        end

        // pi0830: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0830= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0830= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0830= (i + 830) % 2;  // Phase3: 翻转
          end
        end

        // pi0831: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0831= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0831= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0831= (i + 831) % 2;  // Phase3: 翻转
          end
        end

        // pi0832: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0832= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0832= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0832= (i + 832) % 2;  // Phase3: 翻转
          end
        end

        // pi0833: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0833= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0833= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0833= (i + 833) % 2;  // Phase3: 翻转
          end
        end

        // pi0834: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0834= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0834= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0834= (i + 834) % 2;  // Phase3: 翻转
          end
        end

        // pi0835: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0835= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0835= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0835= (i + 835) % 2;  // Phase3: 翻转
          end
        end

        // pi0836: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0836= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0836= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0836= (i + 836) % 2;  // Phase3: 翻转
          end
        end

        // pi0837: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0837= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0837= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0837= (i + 837) % 2;  // Phase3: 翻转
          end
        end

        // pi0838: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0838= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0838= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0838= (i + 838) % 2;  // Phase3: 翻转
          end
        end

        // pi0839: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0839= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0839= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0839= (i + 839) % 2;  // Phase3: 翻转
          end
        end

        // pi0840: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0840= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0840= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0840= (i + 840) % 2;  // Phase3: 翻转
          end
        end

        // pi0841: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0841= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0841= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0841= (i + 841) % 2;  // Phase3: 翻转
          end
        end

        // pi0842: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0842= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0842= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0842= (i + 842) % 2;  // Phase3: 翻转
          end
        end

        // pi0843: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0843= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0843= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0843= (i + 843) % 2;  // Phase3: 翻转
          end
        end

        // pi0844: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0844= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0844= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0844= (i + 844) % 2;  // Phase3: 翻转
          end
        end

        // pi0845: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0845= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0845= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0845= (i + 845) % 2;  // Phase3: 翻转
          end
        end

        // pi0846: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0846= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0846= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0846= (i + 846) % 2;  // Phase3: 翻转
          end
        end

        // pi0847: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0847= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0847= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0847= (i + 847) % 2;  // Phase3: 翻转
          end
        end

        // pi0848: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0848= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0848= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0848= (i + 848) % 2;  // Phase3: 翻转
          end
        end

        // pi0849: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0849= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0849= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0849= (i + 849) % 2;  // Phase3: 翻转
          end
        end

        // pi0850: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0850= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0850= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0850= (i + 850) % 2;  // Phase3: 翻转
          end
        end

        // pi0851: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0851= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0851= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0851= (i + 851) % 2;  // Phase3: 翻转
          end
        end

        // pi0852: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0852= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0852= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0852= (i + 852) % 2;  // Phase3: 翻转
          end
        end

        // pi0853: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0853= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0853= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0853= (i + 853) % 2;  // Phase3: 翻转
          end
        end

        // pi0854: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0854= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0854= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0854= (i + 854) % 2;  // Phase3: 翻转
          end
        end

        // pi0855: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0855= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0855= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0855= (i + 855) % 2;  // Phase3: 翻转
          end
        end

        // pi0856: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0856= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0856= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0856= (i + 856) % 2;  // Phase3: 翻转
          end
        end

        // pi0857: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0857= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0857= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0857= (i + 857) % 2;  // Phase3: 翻转
          end
        end

        // pi0858: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0858= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0858= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0858= (i + 858) % 2;  // Phase3: 翻转
          end
        end

        // pi0859: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0859= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0859= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0859= (i + 859) % 2;  // Phase3: 翻转
          end
        end

        // pi0860: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0860= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0860= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0860= (i + 860) % 2;  // Phase3: 翻转
          end
        end

        // pi0861: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0861= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0861= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0861= (i + 861) % 2;  // Phase3: 翻转
          end
        end

        // pi0862: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0862= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0862= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0862= (i + 862) % 2;  // Phase3: 翻转
          end
        end

        // pi0863: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0863= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0863= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0863= (i + 863) % 2;  // Phase3: 翻转
          end
        end

        // pi0864: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0864= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0864= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0864= (i + 864) % 2;  // Phase3: 翻转
          end
        end

        // pi0865: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0865= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0865= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0865= (i + 865) % 2;  // Phase3: 翻转
          end
        end

        // pi0866: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0866= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0866= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0866= (i + 866) % 2;  // Phase3: 翻转
          end
        end

        // pi0867: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0867= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0867= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0867= (i + 867) % 2;  // Phase3: 翻转
          end
        end

        // pi0868: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0868= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0868= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0868= (i + 868) % 2;  // Phase3: 翻转
          end
        end

        // pi0869: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0869= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0869= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0869= (i + 869) % 2;  // Phase3: 翻转
          end
        end

        // pi0870: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0870= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0870= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0870= (i + 870) % 2;  // Phase3: 翻转
          end
        end

        // pi0871: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0871= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0871= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0871= (i + 871) % 2;  // Phase3: 翻转
          end
        end

        // pi0872: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0872= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0872= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0872= (i + 872) % 2;  // Phase3: 翻转
          end
        end

        // pi0873: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0873= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0873= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0873= (i + 873) % 2;  // Phase3: 翻转
          end
        end

        // pi0874: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0874= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0874= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0874= (i + 874) % 2;  // Phase3: 翻转
          end
        end

        // pi0875: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0875= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0875= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0875= (i + 875) % 2;  // Phase3: 翻转
          end
        end

        // pi0876: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0876= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0876= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0876= (i + 876) % 2;  // Phase3: 翻转
          end
        end

        // pi0877: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0877= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0877= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0877= (i + 877) % 2;  // Phase3: 翻转
          end
        end

        // pi0878: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0878= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0878= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0878= (i + 878) % 2;  // Phase3: 翻转
          end
        end

        // pi0879: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0879= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0879= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0879= (i + 879) % 2;  // Phase3: 翻转
          end
        end

        // pi0880: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0880= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0880= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0880= (i + 880) % 2;  // Phase3: 翻转
          end
        end

        // pi0881: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0881= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0881= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0881= (i + 881) % 2;  // Phase3: 翻转
          end
        end

        // pi0882: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0882= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0882= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0882= (i + 882) % 2;  // Phase3: 翻转
          end
        end

        // pi0883: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0883= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0883= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0883= (i + 883) % 2;  // Phase3: 翻转
          end
        end

        // pi0884: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0884= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0884= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0884= (i + 884) % 2;  // Phase3: 翻转
          end
        end

        // pi0885: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0885= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0885= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0885= (i + 885) % 2;  // Phase3: 翻转
          end
        end

        // pi0886: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0886= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0886= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0886= (i + 886) % 2;  // Phase3: 翻转
          end
        end

        // pi0887: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0887= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0887= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0887= (i + 887) % 2;  // Phase3: 翻转
          end
        end

        // pi0888: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0888= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0888= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0888= (i + 888) % 2;  // Phase3: 翻转
          end
        end

        // pi0889: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0889= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0889= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0889= (i + 889) % 2;  // Phase3: 翻转
          end
        end

        // pi0890: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0890= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0890= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0890= (i + 890) % 2;  // Phase3: 翻转
          end
        end

        // pi0891: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0891= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0891= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0891= (i + 891) % 2;  // Phase3: 翻转
          end
        end

        // pi0892: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0892= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0892= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0892= (i + 892) % 2;  // Phase3: 翻转
          end
        end

        // pi0893: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0893= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0893= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0893= (i + 893) % 2;  // Phase3: 翻转
          end
        end

        // pi0894: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0894= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0894= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0894= (i + 894) % 2;  // Phase3: 翻转
          end
        end

        // pi0895: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0895= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0895= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0895= (i + 895) % 2;  // Phase3: 翻转
          end
        end

        // pi0896: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0896= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0896= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0896= (i + 896) % 2;  // Phase3: 翻转
          end
        end

        // pi0897: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0897= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0897= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0897= (i + 897) % 2;  // Phase3: 翻转
          end
        end

        // pi0898: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0898= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0898= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0898= (i + 898) % 2;  // Phase3: 翻转
          end
        end

        // pi0899: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0899= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0899= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0899= (i + 899) % 2;  // Phase3: 翻转
          end
        end

        // pi0900: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0900= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0900= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0900= (i + 900) % 2;  // Phase3: 翻转
          end
        end

        // pi0901: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0901= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0901= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0901= (i + 901) % 2;  // Phase3: 翻转
          end
        end

        // pi0902: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0902= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0902= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0902= (i + 902) % 2;  // Phase3: 翻转
          end
        end

        // pi0903: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0903= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0903= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0903= (i + 903) % 2;  // Phase3: 翻转
          end
        end

        // pi0904: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0904= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0904= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0904= (i + 904) % 2;  // Phase3: 翻转
          end
        end

        // pi0905: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0905= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0905= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0905= (i + 905) % 2;  // Phase3: 翻转
          end
        end

        // pi0906: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0906= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0906= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0906= (i + 906) % 2;  // Phase3: 翻转
          end
        end

        // pi0907: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0907= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0907= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0907= (i + 907) % 2;  // Phase3: 翻转
          end
        end

        // pi0908: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0908= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0908= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0908= (i + 908) % 2;  // Phase3: 翻转
          end
        end

        // pi0909: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0909= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0909= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0909= (i + 909) % 2;  // Phase3: 翻转
          end
        end

        // pi0910: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0910= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0910= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0910= (i + 910) % 2;  // Phase3: 翻转
          end
        end

        // pi0911: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0911= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0911= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0911= (i + 911) % 2;  // Phase3: 翻转
          end
        end

        // pi0912: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0912= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0912= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0912= (i + 912) % 2;  // Phase3: 翻转
          end
        end

        // pi0913: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0913= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0913= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0913= (i + 913) % 2;  // Phase3: 翻转
          end
        end

        // pi0914: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0914= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0914= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0914= (i + 914) % 2;  // Phase3: 翻转
          end
        end

        // pi0915: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0915= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0915= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0915= (i + 915) % 2;  // Phase3: 翻转
          end
        end

        // pi0916: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0916= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0916= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0916= (i + 916) % 2;  // Phase3: 翻转
          end
        end

        // pi0917: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0917= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0917= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0917= (i + 917) % 2;  // Phase3: 翻转
          end
        end

        // pi0918: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0918= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0918= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0918= (i + 918) % 2;  // Phase3: 翻转
          end
        end

        // pi0919: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0919= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0919= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0919= (i + 919) % 2;  // Phase3: 翻转
          end
        end

        // pi0920: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0920= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0920= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0920= (i + 920) % 2;  // Phase3: 翻转
          end
        end

        // pi0921: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0921= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0921= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0921= (i + 921) % 2;  // Phase3: 翻转
          end
        end

        // pi0922: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0922= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0922= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0922= (i + 922) % 2;  // Phase3: 翻转
          end
        end

        // pi0923: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0923= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0923= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0923= (i + 923) % 2;  // Phase3: 翻转
          end
        end

        // pi0924: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0924= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0924= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0924= (i + 924) % 2;  // Phase3: 翻转
          end
        end

        // pi0925: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0925= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0925= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0925= (i + 925) % 2;  // Phase3: 翻转
          end
        end

        // pi0926: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0926= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0926= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0926= (i + 926) % 2;  // Phase3: 翻转
          end
        end

        // pi0927: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0927= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0927= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0927= (i + 927) % 2;  // Phase3: 翻转
          end
        end

        // pi0928: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0928= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0928= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0928= (i + 928) % 2;  // Phase3: 翻转
          end
        end

        // pi0929: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0929= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0929= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0929= (i + 929) % 2;  // Phase3: 翻转
          end
        end

        // pi0930: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0930= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0930= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0930= (i + 930) % 2;  // Phase3: 翻转
          end
        end

        // pi0931: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0931= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0931= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0931= (i + 931) % 2;  // Phase3: 翻转
          end
        end

        // pi0932: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0932= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0932= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0932= (i + 932) % 2;  // Phase3: 翻转
          end
        end

        // pi0933: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0933= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0933= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0933= (i + 933) % 2;  // Phase3: 翻转
          end
        end

        // pi0934: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0934= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0934= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0934= (i + 934) % 2;  // Phase3: 翻转
          end
        end

        // pi0935: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0935= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0935= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0935= (i + 935) % 2;  // Phase3: 翻转
          end
        end

        // pi0936: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0936= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0936= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0936= (i + 936) % 2;  // Phase3: 翻转
          end
        end

        // pi0937: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0937= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0937= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0937= (i + 937) % 2;  // Phase3: 翻转
          end
        end

        // pi0938: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0938= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0938= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0938= (i + 938) % 2;  // Phase3: 翻转
          end
        end

        // pi0939: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0939= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0939= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0939= (i + 939) % 2;  // Phase3: 翻转
          end
        end

        // pi0940: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0940= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0940= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0940= (i + 940) % 2;  // Phase3: 翻转
          end
        end

        // pi0941: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0941= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0941= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0941= (i + 941) % 2;  // Phase3: 翻转
          end
        end

        // pi0942: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0942= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0942= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0942= (i + 942) % 2;  // Phase3: 翻转
          end
        end

        // pi0943: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0943= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0943= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0943= (i + 943) % 2;  // Phase3: 翻转
          end
        end

        // pi0944: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0944= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0944= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0944= (i + 944) % 2;  // Phase3: 翻转
          end
        end

        // pi0945: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0945= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0945= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0945= (i + 945) % 2;  // Phase3: 翻转
          end
        end

        // pi0946: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0946= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0946= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0946= (i + 946) % 2;  // Phase3: 翻转
          end
        end

        // pi0947: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0947= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0947= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0947= (i + 947) % 2;  // Phase3: 翻转
          end
        end

        // pi0948: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0948= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0948= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0948= (i + 948) % 2;  // Phase3: 翻转
          end
        end

        // pi0949: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0949= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0949= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0949= (i + 949) % 2;  // Phase3: 翻转
          end
        end

        // pi0950: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0950= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0950= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0950= (i + 950) % 2;  // Phase3: 翻转
          end
        end

        // pi0951: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0951= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0951= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0951= (i + 951) % 2;  // Phase3: 翻转
          end
        end

        // pi0952: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0952= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0952= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0952= (i + 952) % 2;  // Phase3: 翻转
          end
        end

        // pi0953: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0953= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0953= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0953= (i + 953) % 2;  // Phase3: 翻转
          end
        end

        // pi0954: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0954= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0954= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0954= (i + 954) % 2;  // Phase3: 翻转
          end
        end

        // pi0955: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0955= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0955= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0955= (i + 955) % 2;  // Phase3: 翻转
          end
        end

        // pi0956: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0956= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0956= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0956= (i + 956) % 2;  // Phase3: 翻转
          end
        end

        // pi0957: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0957= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0957= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0957= (i + 957) % 2;  // Phase3: 翻转
          end
        end

        // pi0958: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0958= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0958= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0958= (i + 958) % 2;  // Phase3: 翻转
          end
        end

        // pi0959: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0959= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0959= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0959= (i + 959) % 2;  // Phase3: 翻转
          end
        end

        // pi0960: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0960= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0960= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0960= (i + 960) % 2;  // Phase3: 翻转
          end
        end

        // pi0961: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0961= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0961= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0961= (i + 961) % 2;  // Phase3: 翻转
          end
        end

        // pi0962: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0962= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0962= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0962= (i + 962) % 2;  // Phase3: 翻转
          end
        end

        // pi0963: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0963= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0963= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0963= (i + 963) % 2;  // Phase3: 翻转
          end
        end

        // pi0964: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0964= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0964= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0964= (i + 964) % 2;  // Phase3: 翻转
          end
        end

        // pi0965: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0965= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0965= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0965= (i + 965) % 2;  // Phase3: 翻转
          end
        end

        // pi0966: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0966= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0966= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0966= (i + 966) % 2;  // Phase3: 翻转
          end
        end

        // pi0967: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0967= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0967= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0967= (i + 967) % 2;  // Phase3: 翻转
          end
        end

        // pi0968: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0968= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0968= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0968= (i + 968) % 2;  // Phase3: 翻转
          end
        end

        // pi0969: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0969= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0969= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0969= (i + 969) % 2;  // Phase3: 翻转
          end
        end

        // pi0970: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0970= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0970= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0970= (i + 970) % 2;  // Phase3: 翻转
          end
        end

        // pi0971: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0971= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0971= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0971= (i + 971) % 2;  // Phase3: 翻转
          end
        end

        // pi0972: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0972= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0972= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0972= (i + 972) % 2;  // Phase3: 翻转
          end
        end

        // pi0973: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0973= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0973= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0973= (i + 973) % 2;  // Phase3: 翻转
          end
        end

        // pi0974: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0974= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0974= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0974= (i + 974) % 2;  // Phase3: 翻转
          end
        end

        // pi0975: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0975= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0975= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0975= (i + 975) % 2;  // Phase3: 翻转
          end
        end

        // pi0976: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0976= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0976= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0976= (i + 976) % 2;  // Phase3: 翻转
          end
        end

        // pi0977: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0977= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0977= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0977= (i + 977) % 2;  // Phase3: 翻转
          end
        end

        // pi0978: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0978= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0978= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0978= (i + 978) % 2;  // Phase3: 翻转
          end
        end

        // pi0979: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0979= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0979= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0979= (i + 979) % 2;  // Phase3: 翻转
          end
        end

        // pi0980: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0980= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0980= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0980= (i + 980) % 2;  // Phase3: 翻转
          end
        end

        // pi0981: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0981= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0981= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0981= (i + 981) % 2;  // Phase3: 翻转
          end
        end

        // pi0982: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0982= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0982= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0982= (i + 982) % 2;  // Phase3: 翻转
          end
        end

        // pi0983: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0983= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0983= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0983= (i + 983) % 2;  // Phase3: 翻转
          end
        end

        // pi0984: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0984= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0984= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0984= (i + 984) % 2;  // Phase3: 翻转
          end
        end

        // pi0985: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0985= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0985= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0985= (i + 985) % 2;  // Phase3: 翻转
          end
        end

        // pi0986: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0986= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0986= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0986= (i + 986) % 2;  // Phase3: 翻转
          end
        end

        // pi0987: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0987= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0987= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0987= (i + 987) % 2;  // Phase3: 翻转
          end
        end

        // pi0988: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0988= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0988= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0988= (i + 988) % 2;  // Phase3: 翻转
          end
        end

        // pi0989: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0989= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0989= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0989= (i + 989) % 2;  // Phase3: 翻转
          end
        end

        // pi0990: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0990= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0990= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0990= (i + 990) % 2;  // Phase3: 翻转
          end
        end

        // pi0991: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0991= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0991= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0991= (i + 991) % 2;  // Phase3: 翻转
          end
        end

        // pi0992: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0992= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0992= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0992= (i + 992) % 2;  // Phase3: 翻转
          end
        end

        // pi0993: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0993= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0993= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0993= (i + 993) % 2;  // Phase3: 翻转
          end
        end

        // pi0994: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0994= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0994= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0994= (i + 994) % 2;  // Phase3: 翻转
          end
        end

        // pi0995: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0995= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0995= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0995= (i + 995) % 2;  // Phase3: 翻转
          end
        end

        // pi0996: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0996= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0996= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0996= (i + 996) % 2;  // Phase3: 翻转
          end
        end

        // pi0997: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0997= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0997= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0997= (i + 997) % 2;  // Phase3: 翻转
          end
        end

        // pi0998: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0998= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0998= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0998= (i + 998) % 2;  // Phase3: 翻转
          end
        end

        // pi0999: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi0999= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi0999= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi0999= (i + 999) % 2;  // Phase3: 翻转
          end
        end

        // pi1000: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1000= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1000= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1000= (i + 1000) % 2;  // Phase3: 翻转
          end
        end

        // pi1001: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1001= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1001= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1001= (i + 1001) % 2;  // Phase3: 翻转
          end
        end

        // pi1002: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1002= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1002= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1002= (i + 1002) % 2;  // Phase3: 翻转
          end
        end

        // pi1003: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1003= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1003= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1003= (i + 1003) % 2;  // Phase3: 翻转
          end
        end

        // pi1004: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1004= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1004= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1004= (i + 1004) % 2;  // Phase3: 翻转
          end
        end

        // pi1005: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1005= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1005= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1005= (i + 1005) % 2;  // Phase3: 翻转
          end
        end

        // pi1006: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1006= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1006= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1006= (i + 1006) % 2;  // Phase3: 翻转
          end
        end

        // pi1007: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1007= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1007= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1007= (i + 1007) % 2;  // Phase3: 翻转
          end
        end

        // pi1008: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1008= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1008= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1008= (i + 1008) % 2;  // Phase3: 翻转
          end
        end

        // pi1009: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1009= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1009= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1009= (i + 1009) % 2;  // Phase3: 翻转
          end
        end

        // pi1010: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1010= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1010= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1010= (i + 1010) % 2;  // Phase3: 翻转
          end
        end

        // pi1011: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1011= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1011= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1011= (i + 1011) % 2;  // Phase3: 翻转
          end
        end

        // pi1012: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1012= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1012= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1012= (i + 1012) % 2;  // Phase3: 翻转
          end
        end

        // pi1013: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1013= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1013= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1013= (i + 1013) % 2;  // Phase3: 翻转
          end
        end

        // pi1014: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1014= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1014= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1014= (i + 1014) % 2;  // Phase3: 翻转
          end
        end

        // pi1015: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1015= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1015= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1015= (i + 1015) % 2;  // Phase3: 翻转
          end
        end

        // pi1016: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1016= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1016= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1016= (i + 1016) % 2;  // Phase3: 翻转
          end
        end

        // pi1017: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1017= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1017= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1017= (i + 1017) % 2;  // Phase3: 翻转
          end
        end

        // pi1018: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1018= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1018= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1018= (i + 1018) % 2;  // Phase3: 翻转
          end
        end

        // pi1019: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1019= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1019= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1019= (i + 1019) % 2;  // Phase3: 翻转
          end
        end

        // pi1020: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1020= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1020= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1020= (i + 1020) % 2;  // Phase3: 翻转
          end
        end

        // pi1021: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1021= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1021= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1021= (i + 1021) % 2;  // Phase3: 翻转
          end
        end

        // pi1022: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1022= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1022= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1022= (i + 1022) % 2;  // Phase3: 翻转
          end
        end

        // pi1023: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1023= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1023= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1023= (i + 1023) % 2;  // Phase3: 翻转
          end
        end

        // pi1024: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1024= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1024= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1024= (i + 1024) % 2;  // Phase3: 翻转
          end
        end

        // pi1025: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1025= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1025= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1025= (i + 1025) % 2;  // Phase3: 翻转
          end
        end

        // pi1026: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1026= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1026= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1026= (i + 1026) % 2;  // Phase3: 翻转
          end
        end

        // pi1027: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1027= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1027= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1027= (i + 1027) % 2;  // Phase3: 翻转
          end
        end

        // pi1028: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1028= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1028= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1028= (i + 1028) % 2;  // Phase3: 翻转
          end
        end

        // pi1029: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1029= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1029= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1029= (i + 1029) % 2;  // Phase3: 翻转
          end
        end

        // pi1030: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1030= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1030= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1030= (i + 1030) % 2;  // Phase3: 翻转
          end
        end

        // pi1031: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1031= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1031= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1031= (i + 1031) % 2;  // Phase3: 翻转
          end
        end

        // pi1032: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1032= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1032= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1032= (i + 1032) % 2;  // Phase3: 翻转
          end
        end

        // pi1033: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1033= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1033= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1033= (i + 1033) % 2;  // Phase3: 翻转
          end
        end

        // pi1034: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1034= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1034= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1034= (i + 1034) % 2;  // Phase3: 翻转
          end
        end

        // pi1035: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1035= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1035= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1035= (i + 1035) % 2;  // Phase3: 翻转
          end
        end

        // pi1036: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1036= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1036= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1036= (i + 1036) % 2;  // Phase3: 翻转
          end
        end

        // pi1037: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1037= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1037= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1037= (i + 1037) % 2;  // Phase3: 翻转
          end
        end

        // pi1038: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1038= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1038= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1038= (i + 1038) % 2;  // Phase3: 翻转
          end
        end

        // pi1039: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1039= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1039= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1039= (i + 1039) % 2;  // Phase3: 翻转
          end
        end

        // pi1040: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1040= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1040= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1040= (i + 1040) % 2;  // Phase3: 翻转
          end
        end

        // pi1041: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1041= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1041= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1041= (i + 1041) % 2;  // Phase3: 翻转
          end
        end

        // pi1042: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1042= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1042= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1042= (i + 1042) % 2;  // Phase3: 翻转
          end
        end

        // pi1043: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1043= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1043= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1043= (i + 1043) % 2;  // Phase3: 翻转
          end
        end

        // pi1044: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1044= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1044= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1044= (i + 1044) % 2;  // Phase3: 翻转
          end
        end

        // pi1045: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1045= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1045= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1045= (i + 1045) % 2;  // Phase3: 翻转
          end
        end

        // pi1046: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1046= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1046= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1046= (i + 1046) % 2;  // Phase3: 翻转
          end
        end

        // pi1047: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1047= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1047= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1047= (i + 1047) % 2;  // Phase3: 翻转
          end
        end

        // pi1048: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1048= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1048= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1048= (i + 1048) % 2;  // Phase3: 翻转
          end
        end

        // pi1049: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1049= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1049= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1049= (i + 1049) % 2;  // Phase3: 翻转
          end
        end

        // pi1050: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1050= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1050= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1050= (i + 1050) % 2;  // Phase3: 翻转
          end
        end

        // pi1051: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1051= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1051= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1051= (i + 1051) % 2;  // Phase3: 翻转
          end
        end

        // pi1052: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1052= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1052= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1052= (i + 1052) % 2;  // Phase3: 翻转
          end
        end

        // pi1053: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1053= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1053= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1053= (i + 1053) % 2;  // Phase3: 翻转
          end
        end

        // pi1054: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1054= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1054= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1054= (i + 1054) % 2;  // Phase3: 翻转
          end
        end

        // pi1055: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1055= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1055= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1055= (i + 1055) % 2;  // Phase3: 翻转
          end
        end

        // pi1056: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1056= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1056= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1056= (i + 1056) % 2;  // Phase3: 翻转
          end
        end

        // pi1057: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1057= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1057= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1057= (i + 1057) % 2;  // Phase3: 翻转
          end
        end

        // pi1058: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1058= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1058= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1058= (i + 1058) % 2;  // Phase3: 翻转
          end
        end

        // pi1059: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1059= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1059= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1059= (i + 1059) % 2;  // Phase3: 翻转
          end
        end

        // pi1060: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1060= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1060= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1060= (i + 1060) % 2;  // Phase3: 翻转
          end
        end

        // pi1061: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1061= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1061= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1061= (i + 1061) % 2;  // Phase3: 翻转
          end
        end

        // pi1062: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1062= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1062= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1062= (i + 1062) % 2;  // Phase3: 翻转
          end
        end

        // pi1063: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1063= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1063= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1063= (i + 1063) % 2;  // Phase3: 翻转
          end
        end

        // pi1064: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1064= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1064= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1064= (i + 1064) % 2;  // Phase3: 翻转
          end
        end

        // pi1065: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1065= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1065= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1065= (i + 1065) % 2;  // Phase3: 翻转
          end
        end

        // pi1066: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1066= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1066= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1066= (i + 1066) % 2;  // Phase3: 翻转
          end
        end

        // pi1067: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1067= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1067= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1067= (i + 1067) % 2;  // Phase3: 翻转
          end
        end

        // pi1068: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1068= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1068= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1068= (i + 1068) % 2;  // Phase3: 翻转
          end
        end

        // pi1069: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1069= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1069= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1069= (i + 1069) % 2;  // Phase3: 翻转
          end
        end

        // pi1070: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1070= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1070= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1070= (i + 1070) % 2;  // Phase3: 翻转
          end
        end

        // pi1071: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1071= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1071= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1071= (i + 1071) % 2;  // Phase3: 翻转
          end
        end

        // pi1072: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1072= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1072= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1072= (i + 1072) % 2;  // Phase3: 翻转
          end
        end

        // pi1073: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1073= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1073= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1073= (i + 1073) % 2;  // Phase3: 翻转
          end
        end

        // pi1074: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1074= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1074= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1074= (i + 1074) % 2;  // Phase3: 翻转
          end
        end

        // pi1075: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1075= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1075= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1075= (i + 1075) % 2;  // Phase3: 翻转
          end
        end

        // pi1076: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1076= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1076= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1076= (i + 1076) % 2;  // Phase3: 翻转
          end
        end

        // pi1077: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1077= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1077= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1077= (i + 1077) % 2;  // Phase3: 翻转
          end
        end

        // pi1078: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1078= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1078= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1078= (i + 1078) % 2;  // Phase3: 翻转
          end
        end

        // pi1079: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1079= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1079= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1079= (i + 1079) % 2;  // Phase3: 翻转
          end
        end

        // pi1080: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1080= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1080= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1080= (i + 1080) % 2;  // Phase3: 翻转
          end
        end

        // pi1081: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1081= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1081= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1081= (i + 1081) % 2;  // Phase3: 翻转
          end
        end

        // pi1082: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1082= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1082= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1082= (i + 1082) % 2;  // Phase3: 翻转
          end
        end

        // pi1083: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1083= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1083= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1083= (i + 1083) % 2;  // Phase3: 翻转
          end
        end

        // pi1084: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1084= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1084= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1084= (i + 1084) % 2;  // Phase3: 翻转
          end
        end

        // pi1085: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1085= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1085= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1085= (i + 1085) % 2;  // Phase3: 翻转
          end
        end

        // pi1086: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1086= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1086= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1086= (i + 1086) % 2;  // Phase3: 翻转
          end
        end

        // pi1087: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1087= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1087= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1087= (i + 1087) % 2;  // Phase3: 翻转
          end
        end

        // pi1088: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1088= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1088= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1088= (i + 1088) % 2;  // Phase3: 翻转
          end
        end

        // pi1089: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1089= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1089= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1089= (i + 1089) % 2;  // Phase3: 翻转
          end
        end

        // pi1090: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1090= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1090= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1090= (i + 1090) % 2;  // Phase3: 翻转
          end
        end

        // pi1091: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1091= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1091= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1091= (i + 1091) % 2;  // Phase3: 翻转
          end
        end

        // pi1092: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1092= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1092= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1092= (i + 1092) % 2;  // Phase3: 翻转
          end
        end

        // pi1093: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1093= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1093= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1093= (i + 1093) % 2;  // Phase3: 翻转
          end
        end

        // pi1094: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1094= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1094= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1094= (i + 1094) % 2;  // Phase3: 翻转
          end
        end

        // pi1095: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1095= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1095= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1095= (i + 1095) % 2;  // Phase3: 翻转
          end
        end

        // pi1096: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1096= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1096= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1096= (i + 1096) % 2;  // Phase3: 翻转
          end
        end

        // pi1097: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1097= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1097= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1097= (i + 1097) % 2;  // Phase3: 翻转
          end
        end

        // pi1098: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1098= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1098= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1098= (i + 1098) % 2;  // Phase3: 翻转
          end
        end

        // pi1099: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1099= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1099= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1099= (i + 1099) % 2;  // Phase3: 翻转
          end
        end

        // pi1100: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1100= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1100= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1100= (i + 1100) % 2;  // Phase3: 翻转
          end
        end

        // pi1101: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1101= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1101= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1101= (i + 1101) % 2;  // Phase3: 翻转
          end
        end

        // pi1102: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1102= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1102= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1102= (i + 1102) % 2;  // Phase3: 翻转
          end
        end

        // pi1103: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1103= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1103= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1103= (i + 1103) % 2;  // Phase3: 翻转
          end
        end

        // pi1104: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1104= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1104= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1104= (i + 1104) % 2;  // Phase3: 翻转
          end
        end

        // pi1105: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1105= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1105= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1105= (i + 1105) % 2;  // Phase3: 翻转
          end
        end

        // pi1106: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1106= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1106= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1106= (i + 1106) % 2;  // Phase3: 翻转
          end
        end

        // pi1107: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1107= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1107= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1107= (i + 1107) % 2;  // Phase3: 翻转
          end
        end

        // pi1108: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1108= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1108= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1108= (i + 1108) % 2;  // Phase3: 翻转
          end
        end

        // pi1109: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1109= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1109= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1109= (i + 1109) % 2;  // Phase3: 翻转
          end
        end

        // pi1110: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1110= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1110= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1110= (i + 1110) % 2;  // Phase3: 翻转
          end
        end

        // pi1111: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1111= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1111= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1111= (i + 1111) % 2;  // Phase3: 翻转
          end
        end

        // pi1112: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1112= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1112= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1112= (i + 1112) % 2;  // Phase3: 翻转
          end
        end

        // pi1113: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1113= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1113= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1113= (i + 1113) % 2;  // Phase3: 翻转
          end
        end

        // pi1114: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1114= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1114= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1114= (i + 1114) % 2;  // Phase3: 翻转
          end
        end

        // pi1115: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1115= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1115= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1115= (i + 1115) % 2;  // Phase3: 翻转
          end
        end

        // pi1116: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1116= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1116= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1116= (i + 1116) % 2;  // Phase3: 翻转
          end
        end

        // pi1117: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1117= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1117= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1117= (i + 1117) % 2;  // Phase3: 翻转
          end
        end

        // pi1118: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1118= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1118= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1118= (i + 1118) % 2;  // Phase3: 翻转
          end
        end

        // pi1119: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1119= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1119= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1119= (i + 1119) % 2;  // Phase3: 翻转
          end
        end

        // pi1120: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1120= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1120= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1120= (i + 1120) % 2;  // Phase3: 翻转
          end
        end

        // pi1121: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1121= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1121= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1121= (i + 1121) % 2;  // Phase3: 翻转
          end
        end

        // pi1122: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1122= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1122= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1122= (i + 1122) % 2;  // Phase3: 翻转
          end
        end

        // pi1123: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1123= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1123= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1123= (i + 1123) % 2;  // Phase3: 翻转
          end
        end

        // pi1124: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1124= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1124= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1124= (i + 1124) % 2;  // Phase3: 翻转
          end
        end

        // pi1125: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1125= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1125= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1125= (i + 1125) % 2;  // Phase3: 翻转
          end
        end

        // pi1126: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1126= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1126= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1126= (i + 1126) % 2;  // Phase3: 翻转
          end
        end

        // pi1127: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1127= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1127= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1127= (i + 1127) % 2;  // Phase3: 翻转
          end
        end

        // pi1128: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1128= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1128= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1128= (i + 1128) % 2;  // Phase3: 翻转
          end
        end

        // pi1129: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1129= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1129= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1129= (i + 1129) % 2;  // Phase3: 翻转
          end
        end

        // pi1130: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1130= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1130= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1130= (i + 1130) % 2;  // Phase3: 翻转
          end
        end

        // pi1131: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1131= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1131= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1131= (i + 1131) % 2;  // Phase3: 翻转
          end
        end

        // pi1132: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1132= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1132= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1132= (i + 1132) % 2;  // Phase3: 翻转
          end
        end

        // pi1133: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1133= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1133= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1133= (i + 1133) % 2;  // Phase3: 翻转
          end
        end

        // pi1134: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1134= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1134= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1134= (i + 1134) % 2;  // Phase3: 翻转
          end
        end

        // pi1135: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1135= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1135= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1135= (i + 1135) % 2;  // Phase3: 翻转
          end
        end

        // pi1136: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1136= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1136= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1136= (i + 1136) % 2;  // Phase3: 翻转
          end
        end

        // pi1137: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1137= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1137= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1137= (i + 1137) % 2;  // Phase3: 翻转
          end
        end

        // pi1138: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1138= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1138= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1138= (i + 1138) % 2;  // Phase3: 翻转
          end
        end

        // pi1139: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1139= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1139= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1139= (i + 1139) % 2;  // Phase3: 翻转
          end
        end

        // pi1140: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1140= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1140= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1140= (i + 1140) % 2;  // Phase3: 翻转
          end
        end

        // pi1141: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1141= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1141= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1141= (i + 1141) % 2;  // Phase3: 翻转
          end
        end

        // pi1142: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1142= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1142= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1142= (i + 1142) % 2;  // Phase3: 翻转
          end
        end

        // pi1143: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1143= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1143= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1143= (i + 1143) % 2;  // Phase3: 翻转
          end
        end

        // pi1144: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1144= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1144= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1144= (i + 1144) % 2;  // Phase3: 翻转
          end
        end

        // pi1145: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1145= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1145= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1145= (i + 1145) % 2;  // Phase3: 翻转
          end
        end

        // pi1146: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1146= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1146= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1146= (i + 1146) % 2;  // Phase3: 翻转
          end
        end

        // pi1147: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1147= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1147= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1147= (i + 1147) % 2;  // Phase3: 翻转
          end
        end

        // pi1148: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1148= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1148= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1148= (i + 1148) % 2;  // Phase3: 翻转
          end
        end

        // pi1149: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1149= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1149= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1149= (i + 1149) % 2;  // Phase3: 翻转
          end
        end

        // pi1150: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1150= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1150= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1150= (i + 1150) % 2;  // Phase3: 翻转
          end
        end

        // pi1151: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1151= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1151= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1151= (i + 1151) % 2;  // Phase3: 翻转
          end
        end

        // pi1152: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1152= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1152= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1152= (i + 1152) % 2;  // Phase3: 翻转
          end
        end

        // pi1153: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1153= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1153= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1153= (i + 1153) % 2;  // Phase3: 翻转
          end
        end

        // pi1154: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1154= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1154= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1154= (i + 1154) % 2;  // Phase3: 翻转
          end
        end

        // pi1155: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1155= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1155= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1155= (i + 1155) % 2;  // Phase3: 翻转
          end
        end

        // pi1156: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1156= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1156= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1156= (i + 1156) % 2;  // Phase3: 翻转
          end
        end

        // pi1157: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1157= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1157= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1157= (i + 1157) % 2;  // Phase3: 翻转
          end
        end

        // pi1158: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1158= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1158= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1158= (i + 1158) % 2;  // Phase3: 翻转
          end
        end

        // pi1159: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1159= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1159= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1159= (i + 1159) % 2;  // Phase3: 翻转
          end
        end

        // pi1160: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1160= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1160= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1160= (i + 1160) % 2;  // Phase3: 翻转
          end
        end

        // pi1161: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1161= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1161= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1161= (i + 1161) % 2;  // Phase3: 翻转
          end
        end

        // pi1162: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1162= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1162= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1162= (i + 1162) % 2;  // Phase3: 翻转
          end
        end

        // pi1163: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1163= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1163= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1163= (i + 1163) % 2;  // Phase3: 翻转
          end
        end

        // pi1164: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1164= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1164= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1164= (i + 1164) % 2;  // Phase3: 翻转
          end
        end

        // pi1165: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1165= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1165= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1165= (i + 1165) % 2;  // Phase3: 翻转
          end
        end

        // pi1166: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1166= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1166= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1166= (i + 1166) % 2;  // Phase3: 翻转
          end
        end

        // pi1167: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1167= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1167= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1167= (i + 1167) % 2;  // Phase3: 翻转
          end
        end

        // pi1168: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1168= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1168= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1168= (i + 1168) % 2;  // Phase3: 翻转
          end
        end

        // pi1169: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1169= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1169= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1169= (i + 1169) % 2;  // Phase3: 翻转
          end
        end

        // pi1170: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1170= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1170= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1170= (i + 1170) % 2;  // Phase3: 翻转
          end
        end

        // pi1171: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1171= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1171= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1171= (i + 1171) % 2;  // Phase3: 翻转
          end
        end

        // pi1172: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1172= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1172= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1172= (i + 1172) % 2;  // Phase3: 翻转
          end
        end

        // pi1173: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1173= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1173= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1173= (i + 1173) % 2;  // Phase3: 翻转
          end
        end

        // pi1174: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1174= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1174= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1174= (i + 1174) % 2;  // Phase3: 翻转
          end
        end

        // pi1175: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1175= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1175= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1175= (i + 1175) % 2;  // Phase3: 翻转
          end
        end

        // pi1176: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1176= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1176= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1176= (i + 1176) % 2;  // Phase3: 翻转
          end
        end

        // pi1177: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1177= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1177= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1177= (i + 1177) % 2;  // Phase3: 翻转
          end
        end

        // pi1178: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1178= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1178= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1178= (i + 1178) % 2;  // Phase3: 翻转
          end
        end

        // pi1179: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1179= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1179= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1179= (i + 1179) % 2;  // Phase3: 翻转
          end
        end

        // pi1180: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1180= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1180= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1180= (i + 1180) % 2;  // Phase3: 翻转
          end
        end

        // pi1181: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1181= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1181= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1181= (i + 1181) % 2;  // Phase3: 翻转
          end
        end

        // pi1182: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1182= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1182= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1182= (i + 1182) % 2;  // Phase3: 翻转
          end
        end

        // pi1183: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1183= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1183= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1183= (i + 1183) % 2;  // Phase3: 翻转
          end
        end

        // pi1184: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1184= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1184= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1184= (i + 1184) % 2;  // Phase3: 翻转
          end
        end

        // pi1185: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1185= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1185= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1185= (i + 1185) % 2;  // Phase3: 翻转
          end
        end

        // pi1186: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1186= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1186= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1186= (i + 1186) % 2;  // Phase3: 翻转
          end
        end

        // pi1187: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1187= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1187= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1187= (i + 1187) % 2;  // Phase3: 翻转
          end
        end

        // pi1188: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1188= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1188= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1188= (i + 1188) % 2;  // Phase3: 翻转
          end
        end

        // pi1189: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1189= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1189= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1189= (i + 1189) % 2;  // Phase3: 翻转
          end
        end

        // pi1190: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1190= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1190= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1190= (i + 1190) % 2;  // Phase3: 翻转
          end
        end

        // pi1191: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1191= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1191= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1191= (i + 1191) % 2;  // Phase3: 翻转
          end
        end

        // pi1192: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1192= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1192= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1192= (i + 1192) % 2;  // Phase3: 翻转
          end
        end

        // pi1193: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1193= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1193= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1193= (i + 1193) % 2;  // Phase3: 翻转
          end
        end

        // pi1194: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1194= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1194= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1194= (i + 1194) % 2;  // Phase3: 翻转
          end
        end

        // pi1195: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1195= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1195= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1195= (i + 1195) % 2;  // Phase3: 翻转
          end
        end

        // pi1196: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1196= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1196= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1196= (i + 1196) % 2;  // Phase3: 翻转
          end
        end

        // pi1197: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1197= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1197= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1197= (i + 1197) % 2;  // Phase3: 翻转
          end
        end

        // pi1198: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1198= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1198= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1198= (i + 1198) % 2;  // Phase3: 翻转
          end
        end

        // pi1199: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1199= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1199= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1199= (i + 1199) % 2;  // Phase3: 翻转
          end
        end

        // pi1200: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1200= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1200= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1200= (i + 1200) % 2;  // Phase3: 翻转
          end
        end

        // pi1201: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1201= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1201= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1201= (i + 1201) % 2;  // Phase3: 翻转
          end
        end

        // pi1202: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1202= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1202= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1202= (i + 1202) % 2;  // Phase3: 翻转
          end
        end

        // pi1203: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi1203= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi1203= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi1203= (i + 1203) % 2;  // Phase3: 翻转
          end
        end

      #10;

      if ((i % PRINT_EVERY) == 0) begin
        $display("o_sum=%06x", {po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230});
      end
    end

    $display("o_sum=%06x [final]", {po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230});
    $finish;
  end

  // VCD output
  reg [510:0] dumpfile_name;
  initial begin
    if (!$value$plusargs("DUMPFILE=%s", dumpfile_name)) begin
      $display("Error: No +DUMPFILE argument");
      $finish;
    end
    $display("Dumping VCD to: %s", dumpfile_name);
    $dumpfile(dumpfile_name);
    $dumpvars(0, tb);
  end

  initial begin
    #1;
    $display("FAULT_INJECTED: check_if_force_took_effect");
  end

endmodule
