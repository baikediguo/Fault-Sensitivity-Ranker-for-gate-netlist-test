`timescale 1ns / 1ps

module tb;

  reg \in0[0] ;
  reg \in0[1] ;
  reg \in0[2] ;
  reg \in0[3] ;
  reg \in0[4] ;
  reg \in0[5] ;
  reg \in0[6] ;
  reg \in0[7] ;
  reg \in0[8] ;
  reg \in0[9] ;
  reg \in0[10] ;
  reg \in0[11] ;
  reg \in0[12] ;
  reg \in0[13] ;
  reg \in0[14] ;
  reg \in0[15] ;
  reg \in0[16] ;
  reg \in0[17] ;
  reg \in0[18] ;
  reg \in0[19] ;
  reg \in0[20] ;
  reg \in0[21] ;
  reg \in0[22] ;
  reg \in0[23] ;
  reg \in0[24] ;
  reg \in0[25] ;
  reg \in0[26] ;
  reg \in0[27] ;
  reg \in0[28] ;
  reg \in0[29] ;
  reg \in0[30] ;
  reg \in0[31] ;
  reg \in0[32] ;
  reg \in0[33] ;
  reg \in0[34] ;
  reg \in0[35] ;
  reg \in0[36] ;
  reg \in0[37] ;
  reg \in0[38] ;
  reg \in0[39] ;
  reg \in0[40] ;
  reg \in0[41] ;
  reg \in0[42] ;
  reg \in0[43] ;
  reg \in0[44] ;
  reg \in0[45] ;
  reg \in0[46] ;
  reg \in0[47] ;
  reg \in0[48] ;
  reg \in0[49] ;
  reg \in0[50] ;
  reg \in0[51] ;
  reg \in0[52] ;
  reg \in0[53] ;
  reg \in0[54] ;
  reg \in0[55] ;
  reg \in0[56] ;
  reg \in0[57] ;
  reg \in0[58] ;
  reg \in0[59] ;
  reg \in0[60] ;
  reg \in0[61] ;
  reg \in0[62] ;
  reg \in0[63] ;
  reg \in0[64] ;
  reg \in0[65] ;
  reg \in0[66] ;
  reg \in0[67] ;
  reg \in0[68] ;
  reg \in0[69] ;
  reg \in0[70] ;
  reg \in0[71] ;
  reg \in0[72] ;
  reg \in0[73] ;
  reg \in0[74] ;
  reg \in0[75] ;
  reg \in0[76] ;
  reg \in0[77] ;
  reg \in0[78] ;
  reg \in0[79] ;
  reg \in0[80] ;
  reg \in0[81] ;
  reg \in0[82] ;
  reg \in0[83] ;
  reg \in0[84] ;
  reg \in0[85] ;
  reg \in0[86] ;
  reg \in0[87] ;
  reg \in0[88] ;
  reg \in0[89] ;
  reg \in0[90] ;
  reg \in0[91] ;
  reg \in0[92] ;
  reg \in0[93] ;
  reg \in0[94] ;
  reg \in0[95] ;
  reg \in0[96] ;
  reg \in0[97] ;
  reg \in0[98] ;
  reg \in0[99] ;
  reg \in0[100] ;
  reg \in0[101] ;
  reg \in0[102] ;
  reg \in0[103] ;
  reg \in0[104] ;
  reg \in0[105] ;
  reg \in0[106] ;
  reg \in0[107] ;
  reg \in0[108] ;
  reg \in0[109] ;
  reg \in0[110] ;
  reg \in0[111] ;
  reg \in0[112] ;
  reg \in0[113] ;
  reg \in0[114] ;
  reg \in0[115] ;
  reg \in0[116] ;
  reg \in0[117] ;
  reg \in0[118] ;
  reg \in0[119] ;
  reg \in0[120] ;
  reg \in0[121] ;
  reg \in0[122] ;
  reg \in0[123] ;
  reg \in0[124] ;
  reg \in0[125] ;
  reg \in0[126] ;
  reg \in0[127] ;
  reg \in1[0] ;
  reg \in1[1] ;
  reg \in1[2] ;
  reg \in1[3] ;
  reg \in1[4] ;
  reg \in1[5] ;
  reg \in1[6] ;
  reg \in1[7] ;
  reg \in1[8] ;
  reg \in1[9] ;
  reg \in1[10] ;
  reg \in1[11] ;
  reg \in1[12] ;
  reg \in1[13] ;
  reg \in1[14] ;
  reg \in1[15] ;
  reg \in1[16] ;
  reg \in1[17] ;
  reg \in1[18] ;
  reg \in1[19] ;
  reg \in1[20] ;
  reg \in1[21] ;
  reg \in1[22] ;
  reg \in1[23] ;
  reg \in1[24] ;
  reg \in1[25] ;
  reg \in1[26] ;
  reg \in1[27] ;
  reg \in1[28] ;
  reg \in1[29] ;
  reg \in1[30] ;
  reg \in1[31] ;
  reg \in1[32] ;
  reg \in1[33] ;
  reg \in1[34] ;
  reg \in1[35] ;
  reg \in1[36] ;
  reg \in1[37] ;
  reg \in1[38] ;
  reg \in1[39] ;
  reg \in1[40] ;
  reg \in1[41] ;
  reg \in1[42] ;
  reg \in1[43] ;
  reg \in1[44] ;
  reg \in1[45] ;
  reg \in1[46] ;
  reg \in1[47] ;
  reg \in1[48] ;
  reg \in1[49] ;
  reg \in1[50] ;
  reg \in1[51] ;
  reg \in1[52] ;
  reg \in1[53] ;
  reg \in1[54] ;
  reg \in1[55] ;
  reg \in1[56] ;
  reg \in1[57] ;
  reg \in1[58] ;
  reg \in1[59] ;
  reg \in1[60] ;
  reg \in1[61] ;
  reg \in1[62] ;
  reg \in1[63] ;
  reg \in1[64] ;
  reg \in1[65] ;
  reg \in1[66] ;
  reg \in1[67] ;
  reg \in1[68] ;
  reg \in1[69] ;
  reg \in1[70] ;
  reg \in1[71] ;
  reg \in1[72] ;
  reg \in1[73] ;
  reg \in1[74] ;
  reg \in1[75] ;
  reg \in1[76] ;
  reg \in1[77] ;
  reg \in1[78] ;
  reg \in1[79] ;
  reg \in1[80] ;
  reg \in1[81] ;
  reg \in1[82] ;
  reg \in1[83] ;
  reg \in1[84] ;
  reg \in1[85] ;
  reg \in1[86] ;
  reg \in1[87] ;
  reg \in1[88] ;
  reg \in1[89] ;
  reg \in1[90] ;
  reg \in1[91] ;
  reg \in1[92] ;
  reg \in1[93] ;
  reg \in1[94] ;
  reg \in1[95] ;
  reg \in1[96] ;
  reg \in1[97] ;
  reg \in1[98] ;
  reg \in1[99] ;
  reg \in1[100] ;
  reg \in1[101] ;
  reg \in1[102] ;
  reg \in1[103] ;
  reg \in1[104] ;
  reg \in1[105] ;
  reg \in1[106] ;
  reg \in1[107] ;
  reg \in1[108] ;
  reg \in1[109] ;
  reg \in1[110] ;
  reg \in1[111] ;
  reg \in1[112] ;
  reg \in1[113] ;
  reg \in1[114] ;
  reg \in1[115] ;
  reg \in1[116] ;
  reg \in1[117] ;
  reg \in1[118] ;
  reg \in1[119] ;
  reg \in1[120] ;
  reg \in1[121] ;
  reg \in1[122] ;
  reg \in1[123] ;
  reg \in1[124] ;
  reg \in1[125] ;
  reg \in1[126] ;
  reg \in1[127] ;
  reg \in2[0] ;
  reg \in2[1] ;
  reg \in2[2] ;
  reg \in2[3] ;
  reg \in2[4] ;
  reg \in2[5] ;
  reg \in2[6] ;
  reg \in2[7] ;
  reg \in2[8] ;
  reg \in2[9] ;
  reg \in2[10] ;
  reg \in2[11] ;
  reg \in2[12] ;
  reg \in2[13] ;
  reg \in2[14] ;
  reg \in2[15] ;
  reg \in2[16] ;
  reg \in2[17] ;
  reg \in2[18] ;
  reg \in2[19] ;
  reg \in2[20] ;
  reg \in2[21] ;
  reg \in2[22] ;
  reg \in2[23] ;
  reg \in2[24] ;
  reg \in2[25] ;
  reg \in2[26] ;
  reg \in2[27] ;
  reg \in2[28] ;
  reg \in2[29] ;
  reg \in2[30] ;
  reg \in2[31] ;
  reg \in2[32] ;
  reg \in2[33] ;
  reg \in2[34] ;
  reg \in2[35] ;
  reg \in2[36] ;
  reg \in2[37] ;
  reg \in2[38] ;
  reg \in2[39] ;
  reg \in2[40] ;
  reg \in2[41] ;
  reg \in2[42] ;
  reg \in2[43] ;
  reg \in2[44] ;
  reg \in2[45] ;
  reg \in2[46] ;
  reg \in2[47] ;
  reg \in2[48] ;
  reg \in2[49] ;
  reg \in2[50] ;
  reg \in2[51] ;
  reg \in2[52] ;
  reg \in2[53] ;
  reg \in2[54] ;
  reg \in2[55] ;
  reg \in2[56] ;
  reg \in2[57] ;
  reg \in2[58] ;
  reg \in2[59] ;
  reg \in2[60] ;
  reg \in2[61] ;
  reg \in2[62] ;
  reg \in2[63] ;
  reg \in2[64] ;
  reg \in2[65] ;
  reg \in2[66] ;
  reg \in2[67] ;
  reg \in2[68] ;
  reg \in2[69] ;
  reg \in2[70] ;
  reg \in2[71] ;
  reg \in2[72] ;
  reg \in2[73] ;
  reg \in2[74] ;
  reg \in2[75] ;
  reg \in2[76] ;
  reg \in2[77] ;
  reg \in2[78] ;
  reg \in2[79] ;
  reg \in2[80] ;
  reg \in2[81] ;
  reg \in2[82] ;
  reg \in2[83] ;
  reg \in2[84] ;
  reg \in2[85] ;
  reg \in2[86] ;
  reg \in2[87] ;
  reg \in2[88] ;
  reg \in2[89] ;
  reg \in2[90] ;
  reg \in2[91] ;
  reg \in2[92] ;
  reg \in2[93] ;
  reg \in2[94] ;
  reg \in2[95] ;
  reg \in2[96] ;
  reg \in2[97] ;
  reg \in2[98] ;
  reg \in2[99] ;
  reg \in2[100] ;
  reg \in2[101] ;
  reg \in2[102] ;
  reg \in2[103] ;
  reg \in2[104] ;
  reg \in2[105] ;
  reg \in2[106] ;
  reg \in2[107] ;
  reg \in2[108] ;
  reg \in2[109] ;
  reg \in2[110] ;
  reg \in2[111] ;
  reg \in2[112] ;
  reg \in2[113] ;
  reg \in2[114] ;
  reg \in2[115] ;
  reg \in2[116] ;
  reg \in2[117] ;
  reg \in2[118] ;
  reg \in2[119] ;
  reg \in2[120] ;
  reg \in2[121] ;
  reg \in2[122] ;
  reg \in2[123] ;
  reg \in2[124] ;
  reg \in2[125] ;
  reg \in2[126] ;
  reg \in2[127] ;
  reg \in3[0] ;
  reg \in3[1] ;
  reg \in3[2] ;
  reg \in3[3] ;
  reg \in3[4] ;
  reg \in3[5] ;
  reg \in3[6] ;
  reg \in3[7] ;
  reg \in3[8] ;
  reg \in3[9] ;
  reg \in3[10] ;
  reg \in3[11] ;
  reg \in3[12] ;
  reg \in3[13] ;
  reg \in3[14] ;
  reg \in3[15] ;
  reg \in3[16] ;
  reg \in3[17] ;
  reg \in3[18] ;
  reg \in3[19] ;
  reg \in3[20] ;
  reg \in3[21] ;
  reg \in3[22] ;
  reg \in3[23] ;
  reg \in3[24] ;
  reg \in3[25] ;
  reg \in3[26] ;
  reg \in3[27] ;
  reg \in3[28] ;
  reg \in3[29] ;
  reg \in3[30] ;
  reg \in3[31] ;
  reg \in3[32] ;
  reg \in3[33] ;
  reg \in3[34] ;
  reg \in3[35] ;
  reg \in3[36] ;
  reg \in3[37] ;
  reg \in3[38] ;
  reg \in3[39] ;
  reg \in3[40] ;
  reg \in3[41] ;
  reg \in3[42] ;
  reg \in3[43] ;
  reg \in3[44] ;
  reg \in3[45] ;
  reg \in3[46] ;
  reg \in3[47] ;
  reg \in3[48] ;
  reg \in3[49] ;
  reg \in3[50] ;
  reg \in3[51] ;
  reg \in3[52] ;
  reg \in3[53] ;
  reg \in3[54] ;
  reg \in3[55] ;
  reg \in3[56] ;
  reg \in3[57] ;
  reg \in3[58] ;
  reg \in3[59] ;
  reg \in3[60] ;
  reg \in3[61] ;
  reg \in3[62] ;
  reg \in3[63] ;
  reg \in3[64] ;
  reg \in3[65] ;
  reg \in3[66] ;
  reg \in3[67] ;
  reg \in3[68] ;
  reg \in3[69] ;
  reg \in3[70] ;
  reg \in3[71] ;
  reg \in3[72] ;
  reg \in3[73] ;
  reg \in3[74] ;
  reg \in3[75] ;
  reg \in3[76] ;
  reg \in3[77] ;
  reg \in3[78] ;
  reg \in3[79] ;
  reg \in3[80] ;
  reg \in3[81] ;
  reg \in3[82] ;
  reg \in3[83] ;
  reg \in3[84] ;
  reg \in3[85] ;
  reg \in3[86] ;
  reg \in3[87] ;
  reg \in3[88] ;
  reg \in3[89] ;
  reg \in3[90] ;
  reg \in3[91] ;
  reg \in3[92] ;
  reg \in3[93] ;
  reg \in3[94] ;
  reg \in3[95] ;
  reg \in3[96] ;
  reg \in3[97] ;
  reg \in3[98] ;
  reg \in3[99] ;
  reg \in3[100] ;
  reg \in3[101] ;
  reg \in3[102] ;
  reg \in3[103] ;
  reg \in3[104] ;
  reg \in3[105] ;
  reg \in3[106] ;
  reg \in3[107] ;
  reg \in3[108] ;
  reg \in3[109] ;
  reg \in3[110] ;
  reg \in3[111] ;
  reg \in3[112] ;
  reg \in3[113] ;
  reg \in3[114] ;
  reg \in3[115] ;
  reg \in3[116] ;
  reg \in3[117] ;
  reg \in3[118] ;
  reg \in3[119] ;
  reg \in3[120] ;
  reg \in3[121] ;
  reg \in3[122] ;
  reg \in3[123] ;
  reg \in3[124] ;
  reg \in3[125] ;
  reg \in3[126] ;
  reg \in3[127] ;
  wire \address[0] ;
  wire \address[1] ;
  wire \result[0] ;
  wire \result[1] ;
  wire \result[2] ;
  wire \result[3] ;
  wire \result[4] ;
  wire \result[5] ;
  wire \result[6] ;
  wire \result[7] ;
  wire \result[8] ;
  wire \result[9] ;
  wire \result[10] ;
  wire \result[11] ;
  wire \result[12] ;
  wire \result[13] ;
  wire \result[14] ;
  wire \result[15] ;
  wire \result[16] ;
  wire \result[17] ;
  wire \result[18] ;
  wire \result[19] ;
  wire \result[20] ;
  wire \result[21] ;
  wire \result[22] ;
  wire \result[23] ;
  wire \result[24] ;
  wire \result[25] ;
  wire \result[26] ;
  wire \result[27] ;
  wire \result[28] ;
  wire \result[29] ;
  wire \result[30] ;
  wire \result[31] ;
  wire \result[32] ;
  wire \result[33] ;
  wire \result[34] ;
  wire \result[35] ;
  wire \result[36] ;
  wire \result[37] ;
  wire \result[38] ;
  wire \result[39] ;
  wire \result[40] ;
  wire \result[41] ;
  wire \result[42] ;
  wire \result[43] ;
  wire \result[44] ;
  wire \result[45] ;
  wire \result[46] ;
  wire \result[47] ;
  wire \result[48] ;
  wire \result[49] ;
  wire \result[50] ;
  wire \result[51] ;
  wire \result[52] ;
  wire \result[53] ;
  wire \result[54] ;
  wire \result[55] ;
  wire \result[56] ;
  wire \result[57] ;
  wire \result[58] ;
  wire \result[59] ;
  wire \result[60] ;
  wire \result[61] ;
  wire \result[62] ;
  wire \result[63] ;
  wire \result[64] ;
  wire \result[65] ;
  wire \result[66] ;
  wire \result[67] ;
  wire \result[68] ;
  wire \result[69] ;
  wire \result[70] ;
  wire \result[71] ;
  wire \result[72] ;
  wire \result[73] ;
  wire \result[74] ;
  wire \result[75] ;
  wire \result[76] ;
  wire \result[77] ;
  wire \result[78] ;
  wire \result[79] ;
  wire \result[80] ;
  wire \result[81] ;
  wire \result[82] ;
  wire \result[83] ;
  wire \result[84] ;
  wire \result[85] ;
  wire \result[86] ;
  wire \result[87] ;
  wire \result[88] ;
  wire \result[89] ;
  wire \result[90] ;
  wire \result[91] ;
  wire \result[92] ;
  wire \result[93] ;
  wire \result[94] ;
  wire \result[95] ;
  wire \result[96] ;
  wire \result[97] ;
  wire \result[98] ;
  wire \result[99] ;
  wire \result[100] ;
  wire \result[101] ;
  wire \result[102] ;
  wire \result[103] ;
  wire \result[104] ;
  wire \result[105] ;
  wire \result[106] ;
  wire \result[107] ;
  wire \result[108] ;
  wire \result[109] ;
  wire \result[110] ;
  wire \result[111] ;
  wire \result[112] ;
  wire \result[113] ;
  wire \result[114] ;
  wire \result[115] ;
  wire \result[116] ;
  wire \result[117] ;
  wire \result[118] ;
  wire \result[119] ;
  wire \result[120] ;
  wire \result[121] ;
  wire \result[122] ;
  wire \result[123] ;
  wire \result[124] ;
  wire \result[125] ;
  wire \result[126] ;
  wire \result[127] ;

  top uut (
    .\in0[0] (\in0[0] ),
    .\in0[1] (\in0[1] ),
    .\in0[2] (\in0[2] ),
    .\in0[3] (\in0[3] ),
    .\in0[4] (\in0[4] ),
    .\in0[5] (\in0[5] ),
    .\in0[6] (\in0[6] ),
    .\in0[7] (\in0[7] ),
    .\in0[8] (\in0[8] ),
    .\in0[9] (\in0[9] ),
    .\in0[10] (\in0[10] ),
    .\in0[11] (\in0[11] ),
    .\in0[12] (\in0[12] ),
    .\in0[13] (\in0[13] ),
    .\in0[14] (\in0[14] ),
    .\in0[15] (\in0[15] ),
    .\in0[16] (\in0[16] ),
    .\in0[17] (\in0[17] ),
    .\in0[18] (\in0[18] ),
    .\in0[19] (\in0[19] ),
    .\in0[20] (\in0[20] ),
    .\in0[21] (\in0[21] ),
    .\in0[22] (\in0[22] ),
    .\in0[23] (\in0[23] ),
    .\in0[24] (\in0[24] ),
    .\in0[25] (\in0[25] ),
    .\in0[26] (\in0[26] ),
    .\in0[27] (\in0[27] ),
    .\in0[28] (\in0[28] ),
    .\in0[29] (\in0[29] ),
    .\in0[30] (\in0[30] ),
    .\in0[31] (\in0[31] ),
    .\in0[32] (\in0[32] ),
    .\in0[33] (\in0[33] ),
    .\in0[34] (\in0[34] ),
    .\in0[35] (\in0[35] ),
    .\in0[36] (\in0[36] ),
    .\in0[37] (\in0[37] ),
    .\in0[38] (\in0[38] ),
    .\in0[39] (\in0[39] ),
    .\in0[40] (\in0[40] ),
    .\in0[41] (\in0[41] ),
    .\in0[42] (\in0[42] ),
    .\in0[43] (\in0[43] ),
    .\in0[44] (\in0[44] ),
    .\in0[45] (\in0[45] ),
    .\in0[46] (\in0[46] ),
    .\in0[47] (\in0[47] ),
    .\in0[48] (\in0[48] ),
    .\in0[49] (\in0[49] ),
    .\in0[50] (\in0[50] ),
    .\in0[51] (\in0[51] ),
    .\in0[52] (\in0[52] ),
    .\in0[53] (\in0[53] ),
    .\in0[54] (\in0[54] ),
    .\in0[55] (\in0[55] ),
    .\in0[56] (\in0[56] ),
    .\in0[57] (\in0[57] ),
    .\in0[58] (\in0[58] ),
    .\in0[59] (\in0[59] ),
    .\in0[60] (\in0[60] ),
    .\in0[61] (\in0[61] ),
    .\in0[62] (\in0[62] ),
    .\in0[63] (\in0[63] ),
    .\in0[64] (\in0[64] ),
    .\in0[65] (\in0[65] ),
    .\in0[66] (\in0[66] ),
    .\in0[67] (\in0[67] ),
    .\in0[68] (\in0[68] ),
    .\in0[69] (\in0[69] ),
    .\in0[70] (\in0[70] ),
    .\in0[71] (\in0[71] ),
    .\in0[72] (\in0[72] ),
    .\in0[73] (\in0[73] ),
    .\in0[74] (\in0[74] ),
    .\in0[75] (\in0[75] ),
    .\in0[76] (\in0[76] ),
    .\in0[77] (\in0[77] ),
    .\in0[78] (\in0[78] ),
    .\in0[79] (\in0[79] ),
    .\in0[80] (\in0[80] ),
    .\in0[81] (\in0[81] ),
    .\in0[82] (\in0[82] ),
    .\in0[83] (\in0[83] ),
    .\in0[84] (\in0[84] ),
    .\in0[85] (\in0[85] ),
    .\in0[86] (\in0[86] ),
    .\in0[87] (\in0[87] ),
    .\in0[88] (\in0[88] ),
    .\in0[89] (\in0[89] ),
    .\in0[90] (\in0[90] ),
    .\in0[91] (\in0[91] ),
    .\in0[92] (\in0[92] ),
    .\in0[93] (\in0[93] ),
    .\in0[94] (\in0[94] ),
    .\in0[95] (\in0[95] ),
    .\in0[96] (\in0[96] ),
    .\in0[97] (\in0[97] ),
    .\in0[98] (\in0[98] ),
    .\in0[99] (\in0[99] ),
    .\in0[100] (\in0[100] ),
    .\in0[101] (\in0[101] ),
    .\in0[102] (\in0[102] ),
    .\in0[103] (\in0[103] ),
    .\in0[104] (\in0[104] ),
    .\in0[105] (\in0[105] ),
    .\in0[106] (\in0[106] ),
    .\in0[107] (\in0[107] ),
    .\in0[108] (\in0[108] ),
    .\in0[109] (\in0[109] ),
    .\in0[110] (\in0[110] ),
    .\in0[111] (\in0[111] ),
    .\in0[112] (\in0[112] ),
    .\in0[113] (\in0[113] ),
    .\in0[114] (\in0[114] ),
    .\in0[115] (\in0[115] ),
    .\in0[116] (\in0[116] ),
    .\in0[117] (\in0[117] ),
    .\in0[118] (\in0[118] ),
    .\in0[119] (\in0[119] ),
    .\in0[120] (\in0[120] ),
    .\in0[121] (\in0[121] ),
    .\in0[122] (\in0[122] ),
    .\in0[123] (\in0[123] ),
    .\in0[124] (\in0[124] ),
    .\in0[125] (\in0[125] ),
    .\in0[126] (\in0[126] ),
    .\in0[127] (\in0[127] ),
    .\in1[0] (\in1[0] ),
    .\in1[1] (\in1[1] ),
    .\in1[2] (\in1[2] ),
    .\in1[3] (\in1[3] ),
    .\in1[4] (\in1[4] ),
    .\in1[5] (\in1[5] ),
    .\in1[6] (\in1[6] ),
    .\in1[7] (\in1[7] ),
    .\in1[8] (\in1[8] ),
    .\in1[9] (\in1[9] ),
    .\in1[10] (\in1[10] ),
    .\in1[11] (\in1[11] ),
    .\in1[12] (\in1[12] ),
    .\in1[13] (\in1[13] ),
    .\in1[14] (\in1[14] ),
    .\in1[15] (\in1[15] ),
    .\in1[16] (\in1[16] ),
    .\in1[17] (\in1[17] ),
    .\in1[18] (\in1[18] ),
    .\in1[19] (\in1[19] ),
    .\in1[20] (\in1[20] ),
    .\in1[21] (\in1[21] ),
    .\in1[22] (\in1[22] ),
    .\in1[23] (\in1[23] ),
    .\in1[24] (\in1[24] ),
    .\in1[25] (\in1[25] ),
    .\in1[26] (\in1[26] ),
    .\in1[27] (\in1[27] ),
    .\in1[28] (\in1[28] ),
    .\in1[29] (\in1[29] ),
    .\in1[30] (\in1[30] ),
    .\in1[31] (\in1[31] ),
    .\in1[32] (\in1[32] ),
    .\in1[33] (\in1[33] ),
    .\in1[34] (\in1[34] ),
    .\in1[35] (\in1[35] ),
    .\in1[36] (\in1[36] ),
    .\in1[37] (\in1[37] ),
    .\in1[38] (\in1[38] ),
    .\in1[39] (\in1[39] ),
    .\in1[40] (\in1[40] ),
    .\in1[41] (\in1[41] ),
    .\in1[42] (\in1[42] ),
    .\in1[43] (\in1[43] ),
    .\in1[44] (\in1[44] ),
    .\in1[45] (\in1[45] ),
    .\in1[46] (\in1[46] ),
    .\in1[47] (\in1[47] ),
    .\in1[48] (\in1[48] ),
    .\in1[49] (\in1[49] ),
    .\in1[50] (\in1[50] ),
    .\in1[51] (\in1[51] ),
    .\in1[52] (\in1[52] ),
    .\in1[53] (\in1[53] ),
    .\in1[54] (\in1[54] ),
    .\in1[55] (\in1[55] ),
    .\in1[56] (\in1[56] ),
    .\in1[57] (\in1[57] ),
    .\in1[58] (\in1[58] ),
    .\in1[59] (\in1[59] ),
    .\in1[60] (\in1[60] ),
    .\in1[61] (\in1[61] ),
    .\in1[62] (\in1[62] ),
    .\in1[63] (\in1[63] ),
    .\in1[64] (\in1[64] ),
    .\in1[65] (\in1[65] ),
    .\in1[66] (\in1[66] ),
    .\in1[67] (\in1[67] ),
    .\in1[68] (\in1[68] ),
    .\in1[69] (\in1[69] ),
    .\in1[70] (\in1[70] ),
    .\in1[71] (\in1[71] ),
    .\in1[72] (\in1[72] ),
    .\in1[73] (\in1[73] ),
    .\in1[74] (\in1[74] ),
    .\in1[75] (\in1[75] ),
    .\in1[76] (\in1[76] ),
    .\in1[77] (\in1[77] ),
    .\in1[78] (\in1[78] ),
    .\in1[79] (\in1[79] ),
    .\in1[80] (\in1[80] ),
    .\in1[81] (\in1[81] ),
    .\in1[82] (\in1[82] ),
    .\in1[83] (\in1[83] ),
    .\in1[84] (\in1[84] ),
    .\in1[85] (\in1[85] ),
    .\in1[86] (\in1[86] ),
    .\in1[87] (\in1[87] ),
    .\in1[88] (\in1[88] ),
    .\in1[89] (\in1[89] ),
    .\in1[90] (\in1[90] ),
    .\in1[91] (\in1[91] ),
    .\in1[92] (\in1[92] ),
    .\in1[93] (\in1[93] ),
    .\in1[94] (\in1[94] ),
    .\in1[95] (\in1[95] ),
    .\in1[96] (\in1[96] ),
    .\in1[97] (\in1[97] ),
    .\in1[98] (\in1[98] ),
    .\in1[99] (\in1[99] ),
    .\in1[100] (\in1[100] ),
    .\in1[101] (\in1[101] ),
    .\in1[102] (\in1[102] ),
    .\in1[103] (\in1[103] ),
    .\in1[104] (\in1[104] ),
    .\in1[105] (\in1[105] ),
    .\in1[106] (\in1[106] ),
    .\in1[107] (\in1[107] ),
    .\in1[108] (\in1[108] ),
    .\in1[109] (\in1[109] ),
    .\in1[110] (\in1[110] ),
    .\in1[111] (\in1[111] ),
    .\in1[112] (\in1[112] ),
    .\in1[113] (\in1[113] ),
    .\in1[114] (\in1[114] ),
    .\in1[115] (\in1[115] ),
    .\in1[116] (\in1[116] ),
    .\in1[117] (\in1[117] ),
    .\in1[118] (\in1[118] ),
    .\in1[119] (\in1[119] ),
    .\in1[120] (\in1[120] ),
    .\in1[121] (\in1[121] ),
    .\in1[122] (\in1[122] ),
    .\in1[123] (\in1[123] ),
    .\in1[124] (\in1[124] ),
    .\in1[125] (\in1[125] ),
    .\in1[126] (\in1[126] ),
    .\in1[127] (\in1[127] ),
    .\in2[0] (\in2[0] ),
    .\in2[1] (\in2[1] ),
    .\in2[2] (\in2[2] ),
    .\in2[3] (\in2[3] ),
    .\in2[4] (\in2[4] ),
    .\in2[5] (\in2[5] ),
    .\in2[6] (\in2[6] ),
    .\in2[7] (\in2[7] ),
    .\in2[8] (\in2[8] ),
    .\in2[9] (\in2[9] ),
    .\in2[10] (\in2[10] ),
    .\in2[11] (\in2[11] ),
    .\in2[12] (\in2[12] ),
    .\in2[13] (\in2[13] ),
    .\in2[14] (\in2[14] ),
    .\in2[15] (\in2[15] ),
    .\in2[16] (\in2[16] ),
    .\in2[17] (\in2[17] ),
    .\in2[18] (\in2[18] ),
    .\in2[19] (\in2[19] ),
    .\in2[20] (\in2[20] ),
    .\in2[21] (\in2[21] ),
    .\in2[22] (\in2[22] ),
    .\in2[23] (\in2[23] ),
    .\in2[24] (\in2[24] ),
    .\in2[25] (\in2[25] ),
    .\in2[26] (\in2[26] ),
    .\in2[27] (\in2[27] ),
    .\in2[28] (\in2[28] ),
    .\in2[29] (\in2[29] ),
    .\in2[30] (\in2[30] ),
    .\in2[31] (\in2[31] ),
    .\in2[32] (\in2[32] ),
    .\in2[33] (\in2[33] ),
    .\in2[34] (\in2[34] ),
    .\in2[35] (\in2[35] ),
    .\in2[36] (\in2[36] ),
    .\in2[37] (\in2[37] ),
    .\in2[38] (\in2[38] ),
    .\in2[39] (\in2[39] ),
    .\in2[40] (\in2[40] ),
    .\in2[41] (\in2[41] ),
    .\in2[42] (\in2[42] ),
    .\in2[43] (\in2[43] ),
    .\in2[44] (\in2[44] ),
    .\in2[45] (\in2[45] ),
    .\in2[46] (\in2[46] ),
    .\in2[47] (\in2[47] ),
    .\in2[48] (\in2[48] ),
    .\in2[49] (\in2[49] ),
    .\in2[50] (\in2[50] ),
    .\in2[51] (\in2[51] ),
    .\in2[52] (\in2[52] ),
    .\in2[53] (\in2[53] ),
    .\in2[54] (\in2[54] ),
    .\in2[55] (\in2[55] ),
    .\in2[56] (\in2[56] ),
    .\in2[57] (\in2[57] ),
    .\in2[58] (\in2[58] ),
    .\in2[59] (\in2[59] ),
    .\in2[60] (\in2[60] ),
    .\in2[61] (\in2[61] ),
    .\in2[62] (\in2[62] ),
    .\in2[63] (\in2[63] ),
    .\in2[64] (\in2[64] ),
    .\in2[65] (\in2[65] ),
    .\in2[66] (\in2[66] ),
    .\in2[67] (\in2[67] ),
    .\in2[68] (\in2[68] ),
    .\in2[69] (\in2[69] ),
    .\in2[70] (\in2[70] ),
    .\in2[71] (\in2[71] ),
    .\in2[72] (\in2[72] ),
    .\in2[73] (\in2[73] ),
    .\in2[74] (\in2[74] ),
    .\in2[75] (\in2[75] ),
    .\in2[76] (\in2[76] ),
    .\in2[77] (\in2[77] ),
    .\in2[78] (\in2[78] ),
    .\in2[79] (\in2[79] ),
    .\in2[80] (\in2[80] ),
    .\in2[81] (\in2[81] ),
    .\in2[82] (\in2[82] ),
    .\in2[83] (\in2[83] ),
    .\in2[84] (\in2[84] ),
    .\in2[85] (\in2[85] ),
    .\in2[86] (\in2[86] ),
    .\in2[87] (\in2[87] ),
    .\in2[88] (\in2[88] ),
    .\in2[89] (\in2[89] ),
    .\in2[90] (\in2[90] ),
    .\in2[91] (\in2[91] ),
    .\in2[92] (\in2[92] ),
    .\in2[93] (\in2[93] ),
    .\in2[94] (\in2[94] ),
    .\in2[95] (\in2[95] ),
    .\in2[96] (\in2[96] ),
    .\in2[97] (\in2[97] ),
    .\in2[98] (\in2[98] ),
    .\in2[99] (\in2[99] ),
    .\in2[100] (\in2[100] ),
    .\in2[101] (\in2[101] ),
    .\in2[102] (\in2[102] ),
    .\in2[103] (\in2[103] ),
    .\in2[104] (\in2[104] ),
    .\in2[105] (\in2[105] ),
    .\in2[106] (\in2[106] ),
    .\in2[107] (\in2[107] ),
    .\in2[108] (\in2[108] ),
    .\in2[109] (\in2[109] ),
    .\in2[110] (\in2[110] ),
    .\in2[111] (\in2[111] ),
    .\in2[112] (\in2[112] ),
    .\in2[113] (\in2[113] ),
    .\in2[114] (\in2[114] ),
    .\in2[115] (\in2[115] ),
    .\in2[116] (\in2[116] ),
    .\in2[117] (\in2[117] ),
    .\in2[118] (\in2[118] ),
    .\in2[119] (\in2[119] ),
    .\in2[120] (\in2[120] ),
    .\in2[121] (\in2[121] ),
    .\in2[122] (\in2[122] ),
    .\in2[123] (\in2[123] ),
    .\in2[124] (\in2[124] ),
    .\in2[125] (\in2[125] ),
    .\in2[126] (\in2[126] ),
    .\in2[127] (\in2[127] ),
    .\in3[0] (\in3[0] ),
    .\in3[1] (\in3[1] ),
    .\in3[2] (\in3[2] ),
    .\in3[3] (\in3[3] ),
    .\in3[4] (\in3[4] ),
    .\in3[5] (\in3[5] ),
    .\in3[6] (\in3[6] ),
    .\in3[7] (\in3[7] ),
    .\in3[8] (\in3[8] ),
    .\in3[9] (\in3[9] ),
    .\in3[10] (\in3[10] ),
    .\in3[11] (\in3[11] ),
    .\in3[12] (\in3[12] ),
    .\in3[13] (\in3[13] ),
    .\in3[14] (\in3[14] ),
    .\in3[15] (\in3[15] ),
    .\in3[16] (\in3[16] ),
    .\in3[17] (\in3[17] ),
    .\in3[18] (\in3[18] ),
    .\in3[19] (\in3[19] ),
    .\in3[20] (\in3[20] ),
    .\in3[21] (\in3[21] ),
    .\in3[22] (\in3[22] ),
    .\in3[23] (\in3[23] ),
    .\in3[24] (\in3[24] ),
    .\in3[25] (\in3[25] ),
    .\in3[26] (\in3[26] ),
    .\in3[27] (\in3[27] ),
    .\in3[28] (\in3[28] ),
    .\in3[29] (\in3[29] ),
    .\in3[30] (\in3[30] ),
    .\in3[31] (\in3[31] ),
    .\in3[32] (\in3[32] ),
    .\in3[33] (\in3[33] ),
    .\in3[34] (\in3[34] ),
    .\in3[35] (\in3[35] ),
    .\in3[36] (\in3[36] ),
    .\in3[37] (\in3[37] ),
    .\in3[38] (\in3[38] ),
    .\in3[39] (\in3[39] ),
    .\in3[40] (\in3[40] ),
    .\in3[41] (\in3[41] ),
    .\in3[42] (\in3[42] ),
    .\in3[43] (\in3[43] ),
    .\in3[44] (\in3[44] ),
    .\in3[45] (\in3[45] ),
    .\in3[46] (\in3[46] ),
    .\in3[47] (\in3[47] ),
    .\in3[48] (\in3[48] ),
    .\in3[49] (\in3[49] ),
    .\in3[50] (\in3[50] ),
    .\in3[51] (\in3[51] ),
    .\in3[52] (\in3[52] ),
    .\in3[53] (\in3[53] ),
    .\in3[54] (\in3[54] ),
    .\in3[55] (\in3[55] ),
    .\in3[56] (\in3[56] ),
    .\in3[57] (\in3[57] ),
    .\in3[58] (\in3[58] ),
    .\in3[59] (\in3[59] ),
    .\in3[60] (\in3[60] ),
    .\in3[61] (\in3[61] ),
    .\in3[62] (\in3[62] ),
    .\in3[63] (\in3[63] ),
    .\in3[64] (\in3[64] ),
    .\in3[65] (\in3[65] ),
    .\in3[66] (\in3[66] ),
    .\in3[67] (\in3[67] ),
    .\in3[68] (\in3[68] ),
    .\in3[69] (\in3[69] ),
    .\in3[70] (\in3[70] ),
    .\in3[71] (\in3[71] ),
    .\in3[72] (\in3[72] ),
    .\in3[73] (\in3[73] ),
    .\in3[74] (\in3[74] ),
    .\in3[75] (\in3[75] ),
    .\in3[76] (\in3[76] ),
    .\in3[77] (\in3[77] ),
    .\in3[78] (\in3[78] ),
    .\in3[79] (\in3[79] ),
    .\in3[80] (\in3[80] ),
    .\in3[81] (\in3[81] ),
    .\in3[82] (\in3[82] ),
    .\in3[83] (\in3[83] ),
    .\in3[84] (\in3[84] ),
    .\in3[85] (\in3[85] ),
    .\in3[86] (\in3[86] ),
    .\in3[87] (\in3[87] ),
    .\in3[88] (\in3[88] ),
    .\in3[89] (\in3[89] ),
    .\in3[90] (\in3[90] ),
    .\in3[91] (\in3[91] ),
    .\in3[92] (\in3[92] ),
    .\in3[93] (\in3[93] ),
    .\in3[94] (\in3[94] ),
    .\in3[95] (\in3[95] ),
    .\in3[96] (\in3[96] ),
    .\in3[97] (\in3[97] ),
    .\in3[98] (\in3[98] ),
    .\in3[99] (\in3[99] ),
    .\in3[100] (\in3[100] ),
    .\in3[101] (\in3[101] ),
    .\in3[102] (\in3[102] ),
    .\in3[103] (\in3[103] ),
    .\in3[104] (\in3[104] ),
    .\in3[105] (\in3[105] ),
    .\in3[106] (\in3[106] ),
    .\in3[107] (\in3[107] ),
    .\in3[108] (\in3[108] ),
    .\in3[109] (\in3[109] ),
    .\in3[110] (\in3[110] ),
    .\in3[111] (\in3[111] ),
    .\in3[112] (\in3[112] ),
    .\in3[113] (\in3[113] ),
    .\in3[114] (\in3[114] ),
    .\in3[115] (\in3[115] ),
    .\in3[116] (\in3[116] ),
    .\in3[117] (\in3[117] ),
    .\in3[118] (\in3[118] ),
    .\in3[119] (\in3[119] ),
    .\in3[120] (\in3[120] ),
    .\in3[121] (\in3[121] ),
    .\in3[122] (\in3[122] ),
    .\in3[123] (\in3[123] ),
    .\in3[124] (\in3[124] ),
    .\in3[125] (\in3[125] ),
    .\in3[126] (\in3[126] ),
    .\in3[127] (\in3[127] ),
    .\address[0] (\address[0] ),
    .\address[1] (\address[1] ),
    .\result[0] (\result[0] ),
    .\result[1] (\result[1] ),
    .\result[2] (\result[2] ),
    .\result[3] (\result[3] ),
    .\result[4] (\result[4] ),
    .\result[5] (\result[5] ),
    .\result[6] (\result[6] ),
    .\result[7] (\result[7] ),
    .\result[8] (\result[8] ),
    .\result[9] (\result[9] ),
    .\result[10] (\result[10] ),
    .\result[11] (\result[11] ),
    .\result[12] (\result[12] ),
    .\result[13] (\result[13] ),
    .\result[14] (\result[14] ),
    .\result[15] (\result[15] ),
    .\result[16] (\result[16] ),
    .\result[17] (\result[17] ),
    .\result[18] (\result[18] ),
    .\result[19] (\result[19] ),
    .\result[20] (\result[20] ),
    .\result[21] (\result[21] ),
    .\result[22] (\result[22] ),
    .\result[23] (\result[23] ),
    .\result[24] (\result[24] ),
    .\result[25] (\result[25] ),
    .\result[26] (\result[26] ),
    .\result[27] (\result[27] ),
    .\result[28] (\result[28] ),
    .\result[29] (\result[29] ),
    .\result[30] (\result[30] ),
    .\result[31] (\result[31] ),
    .\result[32] (\result[32] ),
    .\result[33] (\result[33] ),
    .\result[34] (\result[34] ),
    .\result[35] (\result[35] ),
    .\result[36] (\result[36] ),
    .\result[37] (\result[37] ),
    .\result[38] (\result[38] ),
    .\result[39] (\result[39] ),
    .\result[40] (\result[40] ),
    .\result[41] (\result[41] ),
    .\result[42] (\result[42] ),
    .\result[43] (\result[43] ),
    .\result[44] (\result[44] ),
    .\result[45] (\result[45] ),
    .\result[46] (\result[46] ),
    .\result[47] (\result[47] ),
    .\result[48] (\result[48] ),
    .\result[49] (\result[49] ),
    .\result[50] (\result[50] ),
    .\result[51] (\result[51] ),
    .\result[52] (\result[52] ),
    .\result[53] (\result[53] ),
    .\result[54] (\result[54] ),
    .\result[55] (\result[55] ),
    .\result[56] (\result[56] ),
    .\result[57] (\result[57] ),
    .\result[58] (\result[58] ),
    .\result[59] (\result[59] ),
    .\result[60] (\result[60] ),
    .\result[61] (\result[61] ),
    .\result[62] (\result[62] ),
    .\result[63] (\result[63] ),
    .\result[64] (\result[64] ),
    .\result[65] (\result[65] ),
    .\result[66] (\result[66] ),
    .\result[67] (\result[67] ),
    .\result[68] (\result[68] ),
    .\result[69] (\result[69] ),
    .\result[70] (\result[70] ),
    .\result[71] (\result[71] ),
    .\result[72] (\result[72] ),
    .\result[73] (\result[73] ),
    .\result[74] (\result[74] ),
    .\result[75] (\result[75] ),
    .\result[76] (\result[76] ),
    .\result[77] (\result[77] ),
    .\result[78] (\result[78] ),
    .\result[79] (\result[79] ),
    .\result[80] (\result[80] ),
    .\result[81] (\result[81] ),
    .\result[82] (\result[82] ),
    .\result[83] (\result[83] ),
    .\result[84] (\result[84] ),
    .\result[85] (\result[85] ),
    .\result[86] (\result[86] ),
    .\result[87] (\result[87] ),
    .\result[88] (\result[88] ),
    .\result[89] (\result[89] ),
    .\result[90] (\result[90] ),
    .\result[91] (\result[91] ),
    .\result[92] (\result[92] ),
    .\result[93] (\result[93] ),
    .\result[94] (\result[94] ),
    .\result[95] (\result[95] ),
    .\result[96] (\result[96] ),
    .\result[97] (\result[97] ),
    .\result[98] (\result[98] ),
    .\result[99] (\result[99] ),
    .\result[100] (\result[100] ),
    .\result[101] (\result[101] ),
    .\result[102] (\result[102] ),
    .\result[103] (\result[103] ),
    .\result[104] (\result[104] ),
    .\result[105] (\result[105] ),
    .\result[106] (\result[106] ),
    .\result[107] (\result[107] ),
    .\result[108] (\result[108] ),
    .\result[109] (\result[109] ),
    .\result[110] (\result[110] ),
    .\result[111] (\result[111] ),
    .\result[112] (\result[112] ),
    .\result[113] (\result[113] ),
    .\result[114] (\result[114] ),
    .\result[115] (\result[115] ),
    .\result[116] (\result[116] ),
    .\result[117] (\result[117] ),
    .\result[118] (\result[118] ),
    .\result[119] (\result[119] ),
    .\result[120] (\result[120] ),
    .\result[121] (\result[121] ),
    .\result[122] (\result[122] ),
    .\result[123] (\result[123] ),
    .\result[124] (\result[124] ),
    .\result[125] (\result[125] ),
    .\result[126] (\result[126] ),
    .\result[127] (\result[127] )
  );

  integer i;
  parameter STEPS = 1024;

  initial begin
    \in0[0] = 1'b0;
    \in0[1] = 1'b0;
    \in0[2] = 1'b0;
    \in0[3] = 1'b0;
    \in0[4] = 1'b0;
    \in0[5] = 1'b0;
    \in0[6] = 1'b0;
    \in0[7] = 1'b0;
    \in0[8] = 1'b0;
    \in0[9] = 1'b0;
    \in0[10] = 1'b0;
    \in0[11] = 1'b0;
    \in0[12] = 1'b0;
    \in0[13] = 1'b0;
    \in0[14] = 1'b0;
    \in0[15] = 1'b0;
    \in0[16] = 1'b0;
    \in0[17] = 1'b0;
    \in0[18] = 1'b0;
    \in0[19] = 1'b0;
    \in0[20] = 1'b0;
    \in0[21] = 1'b0;
    \in0[22] = 1'b0;
    \in0[23] = 1'b0;
    \in0[24] = 1'b0;
    \in0[25] = 1'b0;
    \in0[26] = 1'b0;
    \in0[27] = 1'b0;
    \in0[28] = 1'b0;
    \in0[29] = 1'b0;
    \in0[30] = 1'b0;
    \in0[31] = 1'b0;
    \in0[32] = 1'b0;
    \in0[33] = 1'b0;
    \in0[34] = 1'b0;
    \in0[35] = 1'b0;
    \in0[36] = 1'b0;
    \in0[37] = 1'b0;
    \in0[38] = 1'b0;
    \in0[39] = 1'b0;
    \in0[40] = 1'b0;
    \in0[41] = 1'b0;
    \in0[42] = 1'b0;
    \in0[43] = 1'b0;
    \in0[44] = 1'b0;
    \in0[45] = 1'b0;
    \in0[46] = 1'b0;
    \in0[47] = 1'b0;
    \in0[48] = 1'b0;
    \in0[49] = 1'b0;
    \in0[50] = 1'b0;
    \in0[51] = 1'b0;
    \in0[52] = 1'b0;
    \in0[53] = 1'b0;
    \in0[54] = 1'b0;
    \in0[55] = 1'b0;
    \in0[56] = 1'b0;
    \in0[57] = 1'b0;
    \in0[58] = 1'b0;
    \in0[59] = 1'b0;
    \in0[60] = 1'b0;
    \in0[61] = 1'b0;
    \in0[62] = 1'b0;
    \in0[63] = 1'b0;
    \in0[64] = 1'b0;
    \in0[65] = 1'b0;
    \in0[66] = 1'b0;
    \in0[67] = 1'b0;
    \in0[68] = 1'b0;
    \in0[69] = 1'b0;
    \in0[70] = 1'b0;
    \in0[71] = 1'b0;
    \in0[72] = 1'b0;
    \in0[73] = 1'b0;
    \in0[74] = 1'b0;
    \in0[75] = 1'b0;
    \in0[76] = 1'b0;
    \in0[77] = 1'b0;
    \in0[78] = 1'b0;
    \in0[79] = 1'b0;
    \in0[80] = 1'b0;
    \in0[81] = 1'b0;
    \in0[82] = 1'b0;
    \in0[83] = 1'b0;
    \in0[84] = 1'b0;
    \in0[85] = 1'b0;
    \in0[86] = 1'b0;
    \in0[87] = 1'b0;
    \in0[88] = 1'b0;
    \in0[89] = 1'b0;
    \in0[90] = 1'b0;
    \in0[91] = 1'b0;
    \in0[92] = 1'b0;
    \in0[93] = 1'b0;
    \in0[94] = 1'b0;
    \in0[95] = 1'b0;
    \in0[96] = 1'b0;
    \in0[97] = 1'b0;
    \in0[98] = 1'b0;
    \in0[99] = 1'b0;
    \in0[100] = 1'b0;
    \in0[101] = 1'b0;
    \in0[102] = 1'b0;
    \in0[103] = 1'b0;
    \in0[104] = 1'b0;
    \in0[105] = 1'b0;
    \in0[106] = 1'b0;
    \in0[107] = 1'b0;
    \in0[108] = 1'b0;
    \in0[109] = 1'b0;
    \in0[110] = 1'b0;
    \in0[111] = 1'b0;
    \in0[112] = 1'b0;
    \in0[113] = 1'b0;
    \in0[114] = 1'b0;
    \in0[115] = 1'b0;
    \in0[116] = 1'b0;
    \in0[117] = 1'b0;
    \in0[118] = 1'b0;
    \in0[119] = 1'b0;
    \in0[120] = 1'b0;
    \in0[121] = 1'b0;
    \in0[122] = 1'b0;
    \in0[123] = 1'b0;
    \in0[124] = 1'b0;
    \in0[125] = 1'b0;
    \in0[126] = 1'b0;
    \in0[127] = 1'b0;
    \in1[0] = 1'b0;
    \in1[1] = 1'b0;
    \in1[2] = 1'b0;
    \in1[3] = 1'b0;
    \in1[4] = 1'b0;
    \in1[5] = 1'b0;
    \in1[6] = 1'b0;
    \in1[7] = 1'b0;
    \in1[8] = 1'b0;
    \in1[9] = 1'b0;
    \in1[10] = 1'b0;
    \in1[11] = 1'b0;
    \in1[12] = 1'b0;
    \in1[13] = 1'b0;
    \in1[14] = 1'b0;
    \in1[15] = 1'b0;
    \in1[16] = 1'b0;
    \in1[17] = 1'b0;
    \in1[18] = 1'b0;
    \in1[19] = 1'b0;
    \in1[20] = 1'b0;
    \in1[21] = 1'b0;
    \in1[22] = 1'b0;
    \in1[23] = 1'b0;
    \in1[24] = 1'b0;
    \in1[25] = 1'b0;
    \in1[26] = 1'b0;
    \in1[27] = 1'b0;
    \in1[28] = 1'b0;
    \in1[29] = 1'b0;
    \in1[30] = 1'b0;
    \in1[31] = 1'b0;
    \in1[32] = 1'b0;
    \in1[33] = 1'b0;
    \in1[34] = 1'b0;
    \in1[35] = 1'b0;
    \in1[36] = 1'b0;
    \in1[37] = 1'b0;
    \in1[38] = 1'b0;
    \in1[39] = 1'b0;
    \in1[40] = 1'b0;
    \in1[41] = 1'b0;
    \in1[42] = 1'b0;
    \in1[43] = 1'b0;
    \in1[44] = 1'b0;
    \in1[45] = 1'b0;
    \in1[46] = 1'b0;
    \in1[47] = 1'b0;
    \in1[48] = 1'b0;
    \in1[49] = 1'b0;
    \in1[50] = 1'b0;
    \in1[51] = 1'b0;
    \in1[52] = 1'b0;
    \in1[53] = 1'b0;
    \in1[54] = 1'b0;
    \in1[55] = 1'b0;
    \in1[56] = 1'b0;
    \in1[57] = 1'b0;
    \in1[58] = 1'b0;
    \in1[59] = 1'b0;
    \in1[60] = 1'b0;
    \in1[61] = 1'b0;
    \in1[62] = 1'b0;
    \in1[63] = 1'b0;
    \in1[64] = 1'b0;
    \in1[65] = 1'b0;
    \in1[66] = 1'b0;
    \in1[67] = 1'b0;
    \in1[68] = 1'b0;
    \in1[69] = 1'b0;
    \in1[70] = 1'b0;
    \in1[71] = 1'b0;
    \in1[72] = 1'b0;
    \in1[73] = 1'b0;
    \in1[74] = 1'b0;
    \in1[75] = 1'b0;
    \in1[76] = 1'b0;
    \in1[77] = 1'b0;
    \in1[78] = 1'b0;
    \in1[79] = 1'b0;
    \in1[80] = 1'b0;
    \in1[81] = 1'b0;
    \in1[82] = 1'b0;
    \in1[83] = 1'b0;
    \in1[84] = 1'b0;
    \in1[85] = 1'b0;
    \in1[86] = 1'b0;
    \in1[87] = 1'b0;
    \in1[88] = 1'b0;
    \in1[89] = 1'b0;
    \in1[90] = 1'b0;
    \in1[91] = 1'b0;
    \in1[92] = 1'b0;
    \in1[93] = 1'b0;
    \in1[94] = 1'b0;
    \in1[95] = 1'b0;
    \in1[96] = 1'b0;
    \in1[97] = 1'b0;
    \in1[98] = 1'b0;
    \in1[99] = 1'b0;
    \in1[100] = 1'b0;
    \in1[101] = 1'b0;
    \in1[102] = 1'b0;
    \in1[103] = 1'b0;
    \in1[104] = 1'b0;
    \in1[105] = 1'b0;
    \in1[106] = 1'b0;
    \in1[107] = 1'b0;
    \in1[108] = 1'b0;
    \in1[109] = 1'b0;
    \in1[110] = 1'b0;
    \in1[111] = 1'b0;
    \in1[112] = 1'b0;
    \in1[113] = 1'b0;
    \in1[114] = 1'b0;
    \in1[115] = 1'b0;
    \in1[116] = 1'b0;
    \in1[117] = 1'b0;
    \in1[118] = 1'b0;
    \in1[119] = 1'b0;
    \in1[120] = 1'b0;
    \in1[121] = 1'b0;
    \in1[122] = 1'b0;
    \in1[123] = 1'b0;
    \in1[124] = 1'b0;
    \in1[125] = 1'b0;
    \in1[126] = 1'b0;
    \in1[127] = 1'b0;
    \in2[0] = 1'b0;
    \in2[1] = 1'b0;
    \in2[2] = 1'b0;
    \in2[3] = 1'b0;
    \in2[4] = 1'b0;
    \in2[5] = 1'b0;
    \in2[6] = 1'b0;
    \in2[7] = 1'b0;
    \in2[8] = 1'b0;
    \in2[9] = 1'b0;
    \in2[10] = 1'b0;
    \in2[11] = 1'b0;
    \in2[12] = 1'b0;
    \in2[13] = 1'b0;
    \in2[14] = 1'b0;
    \in2[15] = 1'b0;
    \in2[16] = 1'b0;
    \in2[17] = 1'b0;
    \in2[18] = 1'b0;
    \in2[19] = 1'b0;
    \in2[20] = 1'b0;
    \in2[21] = 1'b0;
    \in2[22] = 1'b0;
    \in2[23] = 1'b0;
    \in2[24] = 1'b0;
    \in2[25] = 1'b0;
    \in2[26] = 1'b0;
    \in2[27] = 1'b0;
    \in2[28] = 1'b0;
    \in2[29] = 1'b0;
    \in2[30] = 1'b0;
    \in2[31] = 1'b0;
    \in2[32] = 1'b0;
    \in2[33] = 1'b0;
    \in2[34] = 1'b0;
    \in2[35] = 1'b0;
    \in2[36] = 1'b0;
    \in2[37] = 1'b0;
    \in2[38] = 1'b0;
    \in2[39] = 1'b0;
    \in2[40] = 1'b0;
    \in2[41] = 1'b0;
    \in2[42] = 1'b0;
    \in2[43] = 1'b0;
    \in2[44] = 1'b0;
    \in2[45] = 1'b0;
    \in2[46] = 1'b0;
    \in2[47] = 1'b0;
    \in2[48] = 1'b0;
    \in2[49] = 1'b0;
    \in2[50] = 1'b0;
    \in2[51] = 1'b0;
    \in2[52] = 1'b0;
    \in2[53] = 1'b0;
    \in2[54] = 1'b0;
    \in2[55] = 1'b0;
    \in2[56] = 1'b0;
    \in2[57] = 1'b0;
    \in2[58] = 1'b0;
    \in2[59] = 1'b0;
    \in2[60] = 1'b0;
    \in2[61] = 1'b0;
    \in2[62] = 1'b0;
    \in2[63] = 1'b0;
    \in2[64] = 1'b0;
    \in2[65] = 1'b0;
    \in2[66] = 1'b0;
    \in2[67] = 1'b0;
    \in2[68] = 1'b0;
    \in2[69] = 1'b0;
    \in2[70] = 1'b0;
    \in2[71] = 1'b0;
    \in2[72] = 1'b0;
    \in2[73] = 1'b0;
    \in2[74] = 1'b0;
    \in2[75] = 1'b0;
    \in2[76] = 1'b0;
    \in2[77] = 1'b0;
    \in2[78] = 1'b0;
    \in2[79] = 1'b0;
    \in2[80] = 1'b0;
    \in2[81] = 1'b0;
    \in2[82] = 1'b0;
    \in2[83] = 1'b0;
    \in2[84] = 1'b0;
    \in2[85] = 1'b0;
    \in2[86] = 1'b0;
    \in2[87] = 1'b0;
    \in2[88] = 1'b0;
    \in2[89] = 1'b0;
    \in2[90] = 1'b0;
    \in2[91] = 1'b0;
    \in2[92] = 1'b0;
    \in2[93] = 1'b0;
    \in2[94] = 1'b0;
    \in2[95] = 1'b0;
    \in2[96] = 1'b0;
    \in2[97] = 1'b0;
    \in2[98] = 1'b0;
    \in2[99] = 1'b0;
    \in2[100] = 1'b0;
    \in2[101] = 1'b0;
    \in2[102] = 1'b0;
    \in2[103] = 1'b0;
    \in2[104] = 1'b0;
    \in2[105] = 1'b0;
    \in2[106] = 1'b0;
    \in2[107] = 1'b0;
    \in2[108] = 1'b0;
    \in2[109] = 1'b0;
    \in2[110] = 1'b0;
    \in2[111] = 1'b0;
    \in2[112] = 1'b0;
    \in2[113] = 1'b0;
    \in2[114] = 1'b0;
    \in2[115] = 1'b0;
    \in2[116] = 1'b0;
    \in2[117] = 1'b0;
    \in2[118] = 1'b0;
    \in2[119] = 1'b0;
    \in2[120] = 1'b0;
    \in2[121] = 1'b0;
    \in2[122] = 1'b0;
    \in2[123] = 1'b0;
    \in2[124] = 1'b0;
    \in2[125] = 1'b0;
    \in2[126] = 1'b0;
    \in2[127] = 1'b0;
    \in3[0] = 1'b0;
    \in3[1] = 1'b0;
    \in3[2] = 1'b0;
    \in3[3] = 1'b0;
    \in3[4] = 1'b0;
    \in3[5] = 1'b0;
    \in3[6] = 1'b0;
    \in3[7] = 1'b0;
    \in3[8] = 1'b0;
    \in3[9] = 1'b0;
    \in3[10] = 1'b0;
    \in3[11] = 1'b0;
    \in3[12] = 1'b0;
    \in3[13] = 1'b0;
    \in3[14] = 1'b0;
    \in3[15] = 1'b0;
    \in3[16] = 1'b0;
    \in3[17] = 1'b0;
    \in3[18] = 1'b0;
    \in3[19] = 1'b0;
    \in3[20] = 1'b0;
    \in3[21] = 1'b0;
    \in3[22] = 1'b0;
    \in3[23] = 1'b0;
    \in3[24] = 1'b0;
    \in3[25] = 1'b0;
    \in3[26] = 1'b0;
    \in3[27] = 1'b0;
    \in3[28] = 1'b0;
    \in3[29] = 1'b0;
    \in3[30] = 1'b0;
    \in3[31] = 1'b0;
    \in3[32] = 1'b0;
    \in3[33] = 1'b0;
    \in3[34] = 1'b0;
    \in3[35] = 1'b0;
    \in3[36] = 1'b0;
    \in3[37] = 1'b0;
    \in3[38] = 1'b0;
    \in3[39] = 1'b0;
    \in3[40] = 1'b0;
    \in3[41] = 1'b0;
    \in3[42] = 1'b0;
    \in3[43] = 1'b0;
    \in3[44] = 1'b0;
    \in3[45] = 1'b0;
    \in3[46] = 1'b0;
    \in3[47] = 1'b0;
    \in3[48] = 1'b0;
    \in3[49] = 1'b0;
    \in3[50] = 1'b0;
    \in3[51] = 1'b0;
    \in3[52] = 1'b0;
    \in3[53] = 1'b0;
    \in3[54] = 1'b0;
    \in3[55] = 1'b0;
    \in3[56] = 1'b0;
    \in3[57] = 1'b0;
    \in3[58] = 1'b0;
    \in3[59] = 1'b0;
    \in3[60] = 1'b0;
    \in3[61] = 1'b0;
    \in3[62] = 1'b0;
    \in3[63] = 1'b0;
    \in3[64] = 1'b0;
    \in3[65] = 1'b0;
    \in3[66] = 1'b0;
    \in3[67] = 1'b0;
    \in3[68] = 1'b0;
    \in3[69] = 1'b0;
    \in3[70] = 1'b0;
    \in3[71] = 1'b0;
    \in3[72] = 1'b0;
    \in3[73] = 1'b0;
    \in3[74] = 1'b0;
    \in3[75] = 1'b0;
    \in3[76] = 1'b0;
    \in3[77] = 1'b0;
    \in3[78] = 1'b0;
    \in3[79] = 1'b0;
    \in3[80] = 1'b0;
    \in3[81] = 1'b0;
    \in3[82] = 1'b0;
    \in3[83] = 1'b0;
    \in3[84] = 1'b0;
    \in3[85] = 1'b0;
    \in3[86] = 1'b0;
    \in3[87] = 1'b0;
    \in3[88] = 1'b0;
    \in3[89] = 1'b0;
    \in3[90] = 1'b0;
    \in3[91] = 1'b0;
    \in3[92] = 1'b0;
    \in3[93] = 1'b0;
    \in3[94] = 1'b0;
    \in3[95] = 1'b0;
    \in3[96] = 1'b0;
    \in3[97] = 1'b0;
    \in3[98] = 1'b0;
    \in3[99] = 1'b0;
    \in3[100] = 1'b0;
    \in3[101] = 1'b0;
    \in3[102] = 1'b0;
    \in3[103] = 1'b0;
    \in3[104] = 1'b0;
    \in3[105] = 1'b0;
    \in3[106] = 1'b0;
    \in3[107] = 1'b0;
    \in3[108] = 1'b0;
    \in3[109] = 1'b0;
    \in3[110] = 1'b0;
    \in3[111] = 1'b0;
    \in3[112] = 1'b0;
    \in3[113] = 1'b0;
    \in3[114] = 1'b0;
    \in3[115] = 1'b0;
    \in3[116] = 1'b0;
    \in3[117] = 1'b0;
    \in3[118] = 1'b0;
    \in3[119] = 1'b0;
    \in3[120] = 1'b0;
    \in3[121] = 1'b0;
    \in3[122] = 1'b0;
    \in3[123] = 1'b0;
    \in3[124] = 1'b0;
    \in3[125] = 1'b0;
    \in3[126] = 1'b0;
    \in3[127] = 1'b0;

    #10;

    for (i = 0; i < STEPS; i = i + 1) begin
      \in0[112] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[113] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[114] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[115] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[116] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[117] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[118] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[119] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[120] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[121] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[122] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[123] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[124] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[125] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[126] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in0[127] = ((i < 256) ? ((i % 2) < 1) : (i < 512) ? ((i % 4) < 2) : (i < 768) ? ((i % 8) < 4) : ((i % 16) < 8)) ? 1'b1 : 1'b0;
      \in1[112] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[113] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[114] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[115] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[116] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[117] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[118] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[119] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[120] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[121] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[122] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[123] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[124] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[125] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[126] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in1[127] = ((i < 256) ? ((i % 4) < 2) : (i < 512) ? ((i % 8) < 4) : (i < 768) ? ((i % 16) < 8) : ((i % 2) < 1)) ? 1'b1 : 1'b0;
      \in2[112] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[113] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[114] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[115] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[116] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[117] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[118] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[119] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[120] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[121] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[122] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[123] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[124] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[125] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[126] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in2[127] = ((i < 256) ? ((i % 8) < 4) : (i < 512) ? ((i % 16) < 8) : (i < 768) ? ((i % 2) < 1) : ((i % 4) < 2)) ? 1'b1 : 1'b0;
      \in3[112] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[113] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[114] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[115] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[116] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[117] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[118] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[119] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[120] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[121] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[122] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[123] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[124] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[125] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[126] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      \in3[127] = ((i < 256) ? ((i % 16) < 8) : (i < 512) ? ((i % 2) < 1) : (i < 768) ? ((i % 4) < 2) : ((i % 8) < 4)) ? 1'b1 : 1'b0;
      #10;
      $display("o_sum=%0h", {\result[0] , \result[1] , \result[2] , \result[3] , \result[4] , \result[5] , \result[6] , \result[7] , \result[8] , \result[9] , \result[10] , \result[11] , \result[12] , \result[13] , \result[14] , \result[15] , \result[16] , \result[17] , \result[18] , \result[19] , \result[20] , \result[21] , \result[22] , \result[23] , \result[24] , \result[25] , \result[26] , \result[27] , \result[28] , \result[29] , \result[30] , \result[31] , \result[32] , \result[33] , \result[34] , \result[35] , \result[36] , \result[37] , \result[38] , \result[39] , \result[40] , \result[41] , \result[42] , \result[43] , \result[44] , \result[45] , \result[46] , \result[47] , \result[48] , \result[49] , \result[50] , \result[51] , \result[52] , \result[53] , \result[54] , \result[55] , \result[56] , \result[57] , \result[58] , \result[59] , \result[60] , \result[61] , \result[62] , \result[63] , \result[64] , \result[65] , \result[66] , \result[67] , \result[68] , \result[69] , \result[70] , \result[71] , \result[72] , \result[73] , \result[74] , \result[75] , \result[76] , \result[77] , \result[78] , \result[79] , \result[80] , \result[81] , \result[82] , \result[83] , \result[84] , \result[85] , \result[86] , \result[87] , \result[88] , \result[89] , \result[90] , \result[91] , \result[92] , \result[93] , \result[94] , \result[95] , \result[96] , \result[97] , \result[98] , \result[99] , \result[100] , \result[101] , \result[102] , \result[103] , \result[104] , \result[105] , \result[106] , \result[107] , \result[108] , \result[109] , \result[110] , \result[111] , \result[112] , \result[113] , \result[114] , \result[115] , \result[116] , \result[117] , \result[118] , \result[119] , \result[120] , \result[121] , \result[122] , \result[123] , \result[124] , \result[125] , \result[126] , \result[127] , \address[0] , \address[1] });
    end

    $display("o_sum=%0h [final]", {\result[0] , \result[1] , \result[2] , \result[3] , \result[4] , \result[5] , \result[6] , \result[7] , \result[8] , \result[9] , \result[10] , \result[11] , \result[12] , \result[13] , \result[14] , \result[15] , \result[16] , \result[17] , \result[18] , \result[19] , \result[20] , \result[21] , \result[22] , \result[23] , \result[24] , \result[25] , \result[26] , \result[27] , \result[28] , \result[29] , \result[30] , \result[31] , \result[32] , \result[33] , \result[34] , \result[35] , \result[36] , \result[37] , \result[38] , \result[39] , \result[40] , \result[41] , \result[42] , \result[43] , \result[44] , \result[45] , \result[46] , \result[47] , \result[48] , \result[49] , \result[50] , \result[51] , \result[52] , \result[53] , \result[54] , \result[55] , \result[56] , \result[57] , \result[58] , \result[59] , \result[60] , \result[61] , \result[62] , \result[63] , \result[64] , \result[65] , \result[66] , \result[67] , \result[68] , \result[69] , \result[70] , \result[71] , \result[72] , \result[73] , \result[74] , \result[75] , \result[76] , \result[77] , \result[78] , \result[79] , \result[80] , \result[81] , \result[82] , \result[83] , \result[84] , \result[85] , \result[86] , \result[87] , \result[88] , \result[89] , \result[90] , \result[91] , \result[92] , \result[93] , \result[94] , \result[95] , \result[96] , \result[97] , \result[98] , \result[99] , \result[100] , \result[101] , \result[102] , \result[103] , \result[104] , \result[105] , \result[106] , \result[107] , \result[108] , \result[109] , \result[110] , \result[111] , \result[112] , \result[113] , \result[114] , \result[115] , \result[116] , \result[117] , \result[118] , \result[119] , \result[120] , \result[121] , \result[122] , \result[123] , \result[124] , \result[125] , \result[126] , \result[127] , \address[0] , \address[1] });
    $finish;
  end

endmodule