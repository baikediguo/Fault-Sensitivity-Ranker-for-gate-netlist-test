`timescale 1ns / 1ps

module tb;

  reg pi000;
  reg pi001;
  reg pi002;
  reg pi003;
  reg pi004;
  reg pi005;
  reg pi006;
  reg pi007;
  reg pi008;
  reg pi009;
  reg pi010;
  reg pi011;
  reg pi012;
  reg pi013;
  reg pi014;
  reg pi015;
  reg pi016;
  reg pi017;
  reg pi018;
  reg pi019;
  reg pi020;
  reg pi021;
  reg pi022;
  reg pi023;
  reg pi024;
  reg pi025;
  reg pi026;
  reg pi027;
  reg pi028;
  reg pi029;
  reg pi030;
  reg pi031;
  reg pi032;
  reg pi033;
  reg pi034;
  reg pi035;
  reg pi036;
  reg pi037;
  reg pi038;
  reg pi039;
  reg pi040;
  reg pi041;
  reg pi042;
  reg pi043;
  reg pi044;
  reg pi045;
  reg pi046;
  reg pi047;
  reg pi048;
  reg pi049;
  reg pi050;
  reg pi051;
  reg pi052;
  reg pi053;
  reg pi054;
  reg pi055;
  reg pi056;
  reg pi057;
  reg pi058;
  reg pi059;
  reg pi060;
  reg pi061;
  reg pi062;
  reg pi063;
  reg pi064;
  reg pi065;
  reg pi066;
  reg pi067;
  reg pi068;
  reg pi069;
  reg pi070;
  reg pi071;
  reg pi072;
  reg pi073;
  reg pi074;
  reg pi075;
  reg pi076;
  reg pi077;
  reg pi078;
  reg pi079;
  reg pi080;
  reg pi081;
  reg pi082;
  reg pi083;
  reg pi084;
  reg pi085;
  reg pi086;
  reg pi087;
  reg pi088;
  reg pi089;
  reg pi090;
  reg pi091;
  reg pi092;
  reg pi093;
  reg pi094;
  reg pi095;
  reg pi096;
  reg pi097;
  reg pi098;
  reg pi099;
  reg pi100;
  reg pi101;
  reg pi102;
  reg pi103;
  reg pi104;
  reg pi105;
  reg pi106;
  reg pi107;
  reg pi108;
  reg pi109;
  reg pi110;
  reg pi111;
  reg pi112;
  reg pi113;
  reg pi114;
  reg pi115;
  reg pi116;
  reg pi117;
  reg pi118;
  reg pi119;
  reg pi120;
  reg pi121;
  reg pi122;
  reg pi123;
  reg pi124;
  reg pi125;
  reg pi126;
  reg pi127;
  reg pi128;
  reg pi129;
  reg pi130;
  reg pi131;
  reg pi132;
  reg pi133;
  reg pi134;
  reg pi135;
  reg pi136;
  reg pi137;
  reg pi138;
  reg pi139;
  reg pi140;
  reg pi141;
  reg pi142;
  reg pi143;
  reg pi144;
  reg pi145;
  reg pi146;
  wire po000;
  wire po001;
  wire po002;
  wire po003;
  wire po004;
  wire po005;
  wire po006;
  wire po007;
  wire po008;
  wire po009;
  wire po010;
  wire po011;
  wire po012;
  wire po013;
  wire po014;
  wire po015;
  wire po016;
  wire po017;
  wire po018;
  wire po019;
  wire po020;
  wire po021;
  wire po022;
  wire po023;
  wire po024;
  wire po025;
  wire po026;
  wire po027;
  wire po028;
  wire po029;
  wire po030;
  wire po031;
  wire po032;
  wire po033;
  wire po034;
  wire po035;
  wire po036;
  wire po037;
  wire po038;
  wire po039;
  wire po040;
  wire po041;
  wire po042;
  wire po043;
  wire po044;
  wire po045;
  wire po046;
  wire po047;
  wire po048;
  wire po049;
  wire po050;
  wire po051;
  wire po052;
  wire po053;
  wire po054;
  wire po055;
  wire po056;
  wire po057;
  wire po058;
  wire po059;
  wire po060;
  wire po061;
  wire po062;
  wire po063;
  wire po064;
  wire po065;
  wire po066;
  wire po067;
  wire po068;
  wire po069;
  wire po070;
  wire po071;
  wire po072;
  wire po073;
  wire po074;
  wire po075;
  wire po076;
  wire po077;
  wire po078;
  wire po079;
  wire po080;
  wire po081;
  wire po082;
  wire po083;
  wire po084;
  wire po085;
  wire po086;
  wire po087;
  wire po088;
  wire po089;
  wire po090;
  wire po091;
  wire po092;
  wire po093;
  wire po094;
  wire po095;
  wire po096;
  wire po097;
  wire po098;
  wire po099;
  wire po100;
  wire po101;
  wire po102;
  wire po103;
  wire po104;
  wire po105;
  wire po106;
  wire po107;
  wire po108;
  wire po109;
  wire po110;
  wire po111;
  wire po112;
  wire po113;
  wire po114;
  wire po115;
  wire po116;
  wire po117;
  wire po118;
  wire po119;
  wire po120;
  wire po121;
  wire po122;
  wire po123;
  wire po124;
  wire po125;
  wire po126;
  wire po127;
  wire po128;
  wire po129;
  wire po130;
  wire po131;
  wire po132;
  wire po133;
  wire po134;
  wire po135;
  wire po136;
  wire po137;
  wire po138;
  wire po139;
  wire po140;
  wire po141;

  // DUT (combinational)
  i2c uut (
    .pi000(pi000),
    .pi001(pi001),
    .pi002(pi002),
    .pi003(pi003),
    .pi004(pi004),
    .pi005(pi005),
    .pi006(pi006),
    .pi007(pi007),
    .pi008(pi008),
    .pi009(pi009),
    .pi010(pi010),
    .pi011(pi011),
    .pi012(pi012),
    .pi013(pi013),
    .pi014(pi014),
    .pi015(pi015),
    .pi016(pi016),
    .pi017(pi017),
    .pi018(pi018),
    .pi019(pi019),
    .pi020(pi020),
    .pi021(pi021),
    .pi022(pi022),
    .pi023(pi023),
    .pi024(pi024),
    .pi025(pi025),
    .pi026(pi026),
    .pi027(pi027),
    .pi028(pi028),
    .pi029(pi029),
    .pi030(pi030),
    .pi031(pi031),
    .pi032(pi032),
    .pi033(pi033),
    .pi034(pi034),
    .pi035(pi035),
    .pi036(pi036),
    .pi037(pi037),
    .pi038(pi038),
    .pi039(pi039),
    .pi040(pi040),
    .pi041(pi041),
    .pi042(pi042),
    .pi043(pi043),
    .pi044(pi044),
    .pi045(pi045),
    .pi046(pi046),
    .pi047(pi047),
    .pi048(pi048),
    .pi049(pi049),
    .pi050(pi050),
    .pi051(pi051),
    .pi052(pi052),
    .pi053(pi053),
    .pi054(pi054),
    .pi055(pi055),
    .pi056(pi056),
    .pi057(pi057),
    .pi058(pi058),
    .pi059(pi059),
    .pi060(pi060),
    .pi061(pi061),
    .pi062(pi062),
    .pi063(pi063),
    .pi064(pi064),
    .pi065(pi065),
    .pi066(pi066),
    .pi067(pi067),
    .pi068(pi068),
    .pi069(pi069),
    .pi070(pi070),
    .pi071(pi071),
    .pi072(pi072),
    .pi073(pi073),
    .pi074(pi074),
    .pi075(pi075),
    .pi076(pi076),
    .pi077(pi077),
    .pi078(pi078),
    .pi079(pi079),
    .pi080(pi080),
    .pi081(pi081),
    .pi082(pi082),
    .pi083(pi083),
    .pi084(pi084),
    .pi085(pi085),
    .pi086(pi086),
    .pi087(pi087),
    .pi088(pi088),
    .pi089(pi089),
    .pi090(pi090),
    .pi091(pi091),
    .pi092(pi092),
    .pi093(pi093),
    .pi094(pi094),
    .pi095(pi095),
    .pi096(pi096),
    .pi097(pi097),
    .pi098(pi098),
    .pi099(pi099),
    .pi100(pi100),
    .pi101(pi101),
    .pi102(pi102),
    .pi103(pi103),
    .pi104(pi104),
    .pi105(pi105),
    .pi106(pi106),
    .pi107(pi107),
    .pi108(pi108),
    .pi109(pi109),
    .pi110(pi110),
    .pi111(pi111),
    .pi112(pi112),
    .pi113(pi113),
    .pi114(pi114),
    .pi115(pi115),
    .pi116(pi116),
    .pi117(pi117),
    .pi118(pi118),
    .pi119(pi119),
    .pi120(pi120),
    .pi121(pi121),
    .pi122(pi122),
    .pi123(pi123),
    .pi124(pi124),
    .pi125(pi125),
    .pi126(pi126),
    .pi127(pi127),
    .pi128(pi128),
    .pi129(pi129),
    .pi130(pi130),
    .pi131(pi131),
    .pi132(pi132),
    .pi133(pi133),
    .pi134(pi134),
    .pi135(pi135),
    .pi136(pi136),
    .pi137(pi137),
    .pi138(pi138),
    .pi139(pi139),
    .pi140(pi140),
    .pi141(pi141),
    .pi142(pi142),
    .pi143(pi143),
    .pi144(pi144),
    .pi145(pi145),
    .pi146(pi146),
    .po000(po000),
    .po001(po001),
    .po002(po002),
    .po003(po003),
    .po004(po004),
    .po005(po005),
    .po006(po006),
    .po007(po007),
    .po008(po008),
    .po009(po009),
    .po010(po010),
    .po011(po011),
    .po012(po012),
    .po013(po013),
    .po014(po014),
    .po015(po015),
    .po016(po016),
    .po017(po017),
    .po018(po018),
    .po019(po019),
    .po020(po020),
    .po021(po021),
    .po022(po022),
    .po023(po023),
    .po024(po024),
    .po025(po025),
    .po026(po026),
    .po027(po027),
    .po028(po028),
    .po029(po029),
    .po030(po030),
    .po031(po031),
    .po032(po032),
    .po033(po033),
    .po034(po034),
    .po035(po035),
    .po036(po036),
    .po037(po037),
    .po038(po038),
    .po039(po039),
    .po040(po040),
    .po041(po041),
    .po042(po042),
    .po043(po043),
    .po044(po044),
    .po045(po045),
    .po046(po046),
    .po047(po047),
    .po048(po048),
    .po049(po049),
    .po050(po050),
    .po051(po051),
    .po052(po052),
    .po053(po053),
    .po054(po054),
    .po055(po055),
    .po056(po056),
    .po057(po057),
    .po058(po058),
    .po059(po059),
    .po060(po060),
    .po061(po061),
    .po062(po062),
    .po063(po063),
    .po064(po064),
    .po065(po065),
    .po066(po066),
    .po067(po067),
    .po068(po068),
    .po069(po069),
    .po070(po070),
    .po071(po071),
    .po072(po072),
    .po073(po073),
    .po074(po074),
    .po075(po075),
    .po076(po076),
    .po077(po077),
    .po078(po078),
    .po079(po079),
    .po080(po080),
    .po081(po081),
    .po082(po082),
    .po083(po083),
    .po084(po084),
    .po085(po085),
    .po086(po086),
    .po087(po087),
    .po088(po088),
    .po089(po089),
    .po090(po090),
    .po091(po091),
    .po092(po092),
    .po093(po093),
    .po094(po094),
    .po095(po095),
    .po096(po096),
    .po097(po097),
    .po098(po098),
    .po099(po099),
    .po100(po100),
    .po101(po101),
    .po102(po102),
    .po103(po103),
    .po104(po104),
    .po105(po105),
    .po106(po106),
    .po107(po107),
    .po108(po108),
    .po109(po109),
    .po110(po110),
    .po111(po111),
    .po112(po112),
    .po113(po113),
    .po114(po114),
    .po115(po115),
    .po116(po116),
    .po117(po117),
    .po118(po118),
    .po119(po119),
    .po120(po120),
    .po121(po121),
    .po122(po122),
    .po123(po123),
    .po124(po124),
    .po125(po125),
    .po126(po126),
    .po127(po127),
    .po128(po128),
    .po129(po129),
    .po130(po130),
    .po131(po131),
    .po132(po132),
    .po133(po133),
    .po134(po134),
    .po135(po135),
    .po136(po136),
    .po137(po137),
    .po138(po138),
    .po139(po139),
    .po140(po140),
    .po141(po141)
  );

  // Random function
  integer SEED = 6;
  function [7:0] urand(input integer s);
    urand = $random(s) & 8'hFF;
  endfunction

  // Main stimulus (combinational)
  integer i;
  parameter CYCLES = 512;
  parameter PRINT_EVERY = 1;

  initial begin
    pi000= 0;
    pi001= 0;
    pi002= 0;
    pi003= 0;
    pi004= 0;
    pi005= 0;
    pi006= 0;
    pi007= 0;
    pi008= 0;
    pi009= 0;
    pi010= 0;
    pi011= 0;
    pi012= 0;
    pi013= 0;
    pi014= 0;
    pi015= 0;
    pi016= 0;
    pi017= 0;
    pi018= 0;
    pi019= 0;
    pi020= 0;
    pi021= 0;
    pi022= 0;
    pi023= 0;
    pi024= 0;
    pi025= 0;
    pi026= 0;
    pi027= 0;
    pi028= 0;
    pi029= 0;
    pi030= 0;
    pi031= 0;
    pi032= 0;
    pi033= 0;
    pi034= 0;
    pi035= 0;
    pi036= 0;
    pi037= 0;
    pi038= 0;
    pi039= 0;
    pi040= 0;
    pi041= 0;
    pi042= 0;
    pi043= 0;
    pi044= 0;
    pi045= 0;
    pi046= 0;
    pi047= 0;
    pi048= 0;
    pi049= 0;
    pi050= 0;
    pi051= 0;
    pi052= 0;
    pi053= 0;
    pi054= 0;
    pi055= 0;
    pi056= 0;
    pi057= 0;
    pi058= 0;
    pi059= 0;
    pi060= 0;
    pi061= 0;
    pi062= 0;
    pi063= 0;
    pi064= 0;
    pi065= 0;
    pi066= 0;
    pi067= 0;
    pi068= 0;
    pi069= 0;
    pi070= 0;
    pi071= 0;
    pi072= 0;
    pi073= 0;
    pi074= 0;
    pi075= 0;
    pi076= 0;
    pi077= 0;
    pi078= 0;
    pi079= 0;
    pi080= 0;
    pi081= 0;
    pi082= 0;
    pi083= 0;
    pi084= 0;
    pi085= 0;
    pi086= 0;
    pi087= 0;
    pi088= 0;
    pi089= 0;
    pi090= 0;
    pi091= 0;
    pi092= 0;
    pi093= 0;
    pi094= 0;
    pi095= 0;
    pi096= 0;
    pi097= 0;
    pi098= 0;
    pi099= 0;
    pi100= 0;
    pi101= 0;
    pi102= 0;
    pi103= 0;
    pi104= 0;
    pi105= 0;
    pi106= 0;
    pi107= 0;
    pi108= 0;
    pi109= 0;
    pi110= 0;
    pi111= 0;
    pi112= 0;
    pi113= 0;
    pi114= 0;
    pi115= 0;
    pi116= 0;
    pi117= 0;
    pi118= 0;
    pi119= 0;
    pi120= 0;
    pi121= 0;
    pi122= 0;
    pi123= 0;
    pi124= 0;
    pi125= 0;
    pi126= 0;
    pi127= 0;
    pi128= 0;
    pi129= 0;
    pi130= 0;
    pi131= 0;
    pi132= 0;
    pi133= 0;
    pi134= 0;
    pi135= 0;
    pi136= 0;
    pi137= 0;
    pi138= 0;
    pi139= 0;
    pi140= 0;
    pi141= 0;
    pi142= 0;
    pi143= 0;
    pi144= 0;
    pi145= 0;
    pi146= 0;

    #10;

    for (i = 0; i < CYCLES; i = i + 1) begin
        // pi000: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi000= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi000= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi000= (i + 0) % 2;  // Phase3: 翻转
          end
        end

        // pi001: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi001= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi001= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi001= (i + 1) % 2;  // Phase3: 翻转
          end
        end

        // pi002: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi002= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi002= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi002= (i + 2) % 2;  // Phase3: 翻转
          end
        end

        // pi003: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi003= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi003= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi003= (i + 3) % 2;  // Phase3: 翻转
          end
        end

        // pi004: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi004= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi004= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi004= (i + 4) % 2;  // Phase3: 翻转
          end
        end

        // pi005: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi005= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi005= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi005= (i + 5) % 2;  // Phase3: 翻转
          end
        end

        // pi006: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi006= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi006= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi006= (i + 6) % 2;  // Phase3: 翻转
          end
        end

        // pi007: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi007= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi007= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi007= (i + 7) % 2;  // Phase3: 翻转
          end
        end

        // pi008: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi008= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi008= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi008= (i + 8) % 2;  // Phase3: 翻转
          end
        end

        // pi009: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi009= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi009= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi009= (i + 9) % 2;  // Phase3: 翻转
          end
        end

        // pi010: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi010= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi010= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi010= (i + 10) % 2;  // Phase3: 翻转
          end
        end

        // pi011: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi011= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi011= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi011= (i + 11) % 2;  // Phase3: 翻转
          end
        end

        // pi012: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi012= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi012= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi012= (i + 12) % 2;  // Phase3: 翻转
          end
        end

        // pi013: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi013= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi013= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi013= (i + 13) % 2;  // Phase3: 翻转
          end
        end

        // pi014: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi014= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi014= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi014= (i + 14) % 2;  // Phase3: 翻转
          end
        end

        // pi015: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi015= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi015= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi015= (i + 15) % 2;  // Phase3: 翻转
          end
        end

        // pi016: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi016= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi016= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi016= (i + 16) % 2;  // Phase3: 翻转
          end
        end

        // pi017: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi017= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi017= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi017= (i + 17) % 2;  // Phase3: 翻转
          end
        end

        // pi018: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi018= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi018= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi018= (i + 18) % 2;  // Phase3: 翻转
          end
        end

        // pi019: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi019= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi019= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi019= (i + 19) % 2;  // Phase3: 翻转
          end
        end

        // pi020: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi020= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi020= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi020= (i + 20) % 2;  // Phase3: 翻转
          end
        end

        // pi021: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi021= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi021= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi021= (i + 21) % 2;  // Phase3: 翻转
          end
        end

        // pi022: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi022= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi022= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi022= (i + 22) % 2;  // Phase3: 翻转
          end
        end

        // pi023: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi023= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi023= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi023= (i + 23) % 2;  // Phase3: 翻转
          end
        end

        // pi024: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi024= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi024= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi024= (i + 24) % 2;  // Phase3: 翻转
          end
        end

        // pi025: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi025= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi025= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi025= (i + 25) % 2;  // Phase3: 翻转
          end
        end

        // pi026: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi026= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi026= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi026= (i + 26) % 2;  // Phase3: 翻转
          end
        end

        // pi027: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi027= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi027= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi027= (i + 27) % 2;  // Phase3: 翻转
          end
        end

        // pi028: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi028= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi028= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi028= (i + 28) % 2;  // Phase3: 翻转
          end
        end

        // pi029: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi029= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi029= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi029= (i + 29) % 2;  // Phase3: 翻转
          end
        end

        // pi030: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi030= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi030= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi030= (i + 30) % 2;  // Phase3: 翻转
          end
        end

        // pi031: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi031= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi031= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi031= (i + 31) % 2;  // Phase3: 翻转
          end
        end

        // pi032: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi032= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi032= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi032= (i + 32) % 2;  // Phase3: 翻转
          end
        end

        // pi033: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi033= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi033= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi033= (i + 33) % 2;  // Phase3: 翻转
          end
        end

        // pi034: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi034= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi034= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi034= (i + 34) % 2;  // Phase3: 翻转
          end
        end

        // pi035: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi035= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi035= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi035= (i + 35) % 2;  // Phase3: 翻转
          end
        end

        // pi036: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi036= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi036= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi036= (i + 36) % 2;  // Phase3: 翻转
          end
        end

        // pi037: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi037= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi037= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi037= (i + 37) % 2;  // Phase3: 翻转
          end
        end

        // pi038: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi038= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi038= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi038= (i + 38) % 2;  // Phase3: 翻转
          end
        end

        // pi039: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi039= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi039= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi039= (i + 39) % 2;  // Phase3: 翻转
          end
        end

        // pi040: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi040= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi040= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi040= (i + 40) % 2;  // Phase3: 翻转
          end
        end

        // pi041: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi041= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi041= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi041= (i + 41) % 2;  // Phase3: 翻转
          end
        end

        // pi042: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi042= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi042= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi042= (i + 42) % 2;  // Phase3: 翻转
          end
        end

        // pi043: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi043= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi043= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi043= (i + 43) % 2;  // Phase3: 翻转
          end
        end

        // pi044: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi044= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi044= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi044= (i + 44) % 2;  // Phase3: 翻转
          end
        end

        // pi045: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi045= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi045= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi045= (i + 45) % 2;  // Phase3: 翻转
          end
        end

        // pi046: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi046= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi046= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi046= (i + 46) % 2;  // Phase3: 翻转
          end
        end

        // pi047: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi047= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi047= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi047= (i + 47) % 2;  // Phase3: 翻转
          end
        end

        // pi048: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi048= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi048= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi048= (i + 48) % 2;  // Phase3: 翻转
          end
        end

        // pi049: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi049= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi049= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi049= (i + 49) % 2;  // Phase3: 翻转
          end
        end

        // pi050: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi050= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi050= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi050= (i + 50) % 2;  // Phase3: 翻转
          end
        end

        // pi051: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi051= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi051= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi051= (i + 51) % 2;  // Phase3: 翻转
          end
        end

        // pi052: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi052= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi052= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi052= (i + 52) % 2;  // Phase3: 翻转
          end
        end

        // pi053: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi053= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi053= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi053= (i + 53) % 2;  // Phase3: 翻转
          end
        end

        // pi054: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi054= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi054= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi054= (i + 54) % 2;  // Phase3: 翻转
          end
        end

        // pi055: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi055= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi055= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi055= (i + 55) % 2;  // Phase3: 翻转
          end
        end

        // pi056: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi056= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi056= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi056= (i + 56) % 2;  // Phase3: 翻转
          end
        end

        // pi057: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi057= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi057= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi057= (i + 57) % 2;  // Phase3: 翻转
          end
        end

        // pi058: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi058= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi058= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi058= (i + 58) % 2;  // Phase3: 翻转
          end
        end

        // pi059: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi059= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi059= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi059= (i + 59) % 2;  // Phase3: 翻转
          end
        end

        // pi060: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi060= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi060= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi060= (i + 60) % 2;  // Phase3: 翻转
          end
        end

        // pi061: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi061= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi061= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi061= (i + 61) % 2;  // Phase3: 翻转
          end
        end

        // pi062: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi062= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi062= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi062= (i + 62) % 2;  // Phase3: 翻转
          end
        end

        // pi063: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi063= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi063= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi063= (i + 63) % 2;  // Phase3: 翻转
          end
        end

        // pi064: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi064= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi064= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi064= (i + 64) % 2;  // Phase3: 翻转
          end
        end

        // pi065: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi065= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi065= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi065= (i + 65) % 2;  // Phase3: 翻转
          end
        end

        // pi066: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi066= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi066= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi066= (i + 66) % 2;  // Phase3: 翻转
          end
        end

        // pi067: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi067= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi067= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi067= (i + 67) % 2;  // Phase3: 翻转
          end
        end

        // pi068: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi068= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi068= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi068= (i + 68) % 2;  // Phase3: 翻转
          end
        end

        // pi069: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi069= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi069= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi069= (i + 69) % 2;  // Phase3: 翻转
          end
        end

        // pi070: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi070= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi070= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi070= (i + 70) % 2;  // Phase3: 翻转
          end
        end

        // pi071: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi071= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi071= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi071= (i + 71) % 2;  // Phase3: 翻转
          end
        end

        // pi072: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi072= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi072= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi072= (i + 72) % 2;  // Phase3: 翻转
          end
        end

        // pi073: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi073= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi073= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi073= (i + 73) % 2;  // Phase3: 翻转
          end
        end

        // pi074: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi074= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi074= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi074= (i + 74) % 2;  // Phase3: 翻转
          end
        end

        // pi075: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi075= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi075= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi075= (i + 75) % 2;  // Phase3: 翻转
          end
        end

        // pi076: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi076= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi076= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi076= (i + 76) % 2;  // Phase3: 翻转
          end
        end

        // pi077: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi077= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi077= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi077= (i + 77) % 2;  // Phase3: 翻转
          end
        end

        // pi078: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi078= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi078= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi078= (i + 78) % 2;  // Phase3: 翻转
          end
        end

        // pi079: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi079= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi079= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi079= (i + 79) % 2;  // Phase3: 翻转
          end
        end

        // pi080: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi080= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi080= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi080= (i + 80) % 2;  // Phase3: 翻转
          end
        end

        // pi081: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi081= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi081= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi081= (i + 81) % 2;  // Phase3: 翻转
          end
        end

        // pi082: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi082= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi082= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi082= (i + 82) % 2;  // Phase3: 翻转
          end
        end

        // pi083: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi083= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi083= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi083= (i + 83) % 2;  // Phase3: 翻转
          end
        end

        // pi084: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi084= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi084= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi084= (i + 84) % 2;  // Phase3: 翻转
          end
        end

        // pi085: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi085= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi085= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi085= (i + 85) % 2;  // Phase3: 翻转
          end
        end

        // pi086: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi086= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi086= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi086= (i + 86) % 2;  // Phase3: 翻转
          end
        end

        // pi087: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi087= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi087= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi087= (i + 87) % 2;  // Phase3: 翻转
          end
        end

        // pi088: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi088= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi088= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi088= (i + 88) % 2;  // Phase3: 翻转
          end
        end

        // pi089: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi089= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi089= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi089= (i + 89) % 2;  // Phase3: 翻转
          end
        end

        // pi090: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi090= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi090= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi090= (i + 90) % 2;  // Phase3: 翻转
          end
        end

        // pi091: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi091= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi091= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi091= (i + 91) % 2;  // Phase3: 翻转
          end
        end

        // pi092: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi092= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi092= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi092= (i + 92) % 2;  // Phase3: 翻转
          end
        end

        // pi093: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi093= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi093= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi093= (i + 93) % 2;  // Phase3: 翻转
          end
        end

        // pi094: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi094= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi094= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi094= (i + 94) % 2;  // Phase3: 翻转
          end
        end

        // pi095: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi095= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi095= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi095= (i + 95) % 2;  // Phase3: 翻转
          end
        end

        // pi096: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi096= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi096= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi096= (i + 96) % 2;  // Phase3: 翻转
          end
        end

        // pi097: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi097= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi097= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi097= (i + 97) % 2;  // Phase3: 翻转
          end
        end

        // pi098: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi098= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi098= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi098= (i + 98) % 2;  // Phase3: 翻转
          end
        end

        // pi099: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi099= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi099= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi099= (i + 99) % 2;  // Phase3: 翻转
          end
        end

        // pi100: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi100= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi100= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi100= (i + 100) % 2;  // Phase3: 翻转
          end
        end

        // pi101: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi101= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi101= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi101= (i + 101) % 2;  // Phase3: 翻转
          end
        end

        // pi102: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi102= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi102= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi102= (i + 102) % 2;  // Phase3: 翻转
          end
        end

        // pi103: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi103= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi103= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi103= (i + 103) % 2;  // Phase3: 翻转
          end
        end

        // pi104: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi104= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi104= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi104= (i + 104) % 2;  // Phase3: 翻转
          end
        end

        // pi105: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi105= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi105= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi105= (i + 105) % 2;  // Phase3: 翻转
          end
        end

        // pi106: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi106= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi106= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi106= (i + 106) % 2;  // Phase3: 翻转
          end
        end

        // pi107: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi107= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi107= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi107= (i + 107) % 2;  // Phase3: 翻转
          end
        end

        // pi108: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi108= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi108= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi108= (i + 108) % 2;  // Phase3: 翻转
          end
        end

        // pi109: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi109= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi109= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi109= (i + 109) % 2;  // Phase3: 翻转
          end
        end

        // pi110: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi110= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi110= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi110= (i + 110) % 2;  // Phase3: 翻转
          end
        end

        // pi111: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi111= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi111= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi111= (i + 111) % 2;  // Phase3: 翻转
          end
        end

        // pi112: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi112= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi112= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi112= (i + 112) % 2;  // Phase3: 翻转
          end
        end

        // pi113: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi113= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi113= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi113= (i + 113) % 2;  // Phase3: 翻转
          end
        end

        // pi114: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi114= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi114= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi114= (i + 114) % 2;  // Phase3: 翻转
          end
        end

        // pi115: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi115= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi115= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi115= (i + 115) % 2;  // Phase3: 翻转
          end
        end

        // pi116: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi116= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi116= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi116= (i + 116) % 2;  // Phase3: 翻转
          end
        end

        // pi117: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi117= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi117= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi117= (i + 117) % 2;  // Phase3: 翻转
          end
        end

        // pi118: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi118= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi118= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi118= (i + 118) % 2;  // Phase3: 翻转
          end
        end

        // pi119: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi119= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi119= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi119= (i + 119) % 2;  // Phase3: 翻转
          end
        end

        // pi120: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi120= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi120= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi120= (i + 120) % 2;  // Phase3: 翻转
          end
        end

        // pi121: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi121= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi121= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi121= (i + 121) % 2;  // Phase3: 翻转
          end
        end

        // pi122: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi122= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi122= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi122= (i + 122) % 2;  // Phase3: 翻转
          end
        end

        // pi123: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi123= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi123= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi123= (i + 123) % 2;  // Phase3: 翻转
          end
        end

        // pi124: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi124= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi124= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi124= (i + 124) % 2;  // Phase3: 翻转
          end
        end

        // pi125: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi125= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi125= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi125= (i + 125) % 2;  // Phase3: 翻转
          end
        end

        // pi126: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi126= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi126= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi126= (i + 126) % 2;  // Phase3: 翻转
          end
        end

        // pi127: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi127= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi127= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi127= (i + 127) % 2;  // Phase3: 翻转
          end
        end

        // pi128: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi128= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi128= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi128= (i + 128) % 2;  // Phase3: 翻转
          end
        end

        // pi129: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi129= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi129= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi129= (i + 129) % 2;  // Phase3: 翻转
          end
        end

        // pi130: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi130= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi130= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi130= (i + 130) % 2;  // Phase3: 翻转
          end
        end

        // pi131: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi131= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi131= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi131= (i + 131) % 2;  // Phase3: 翻转
          end
        end

        // pi132: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi132= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi132= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi132= (i + 132) % 2;  // Phase3: 翻转
          end
        end

        // pi133: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi133= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi133= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi133= (i + 133) % 2;  // Phase3: 翻转
          end
        end

        // pi134: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi134= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi134= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi134= (i + 134) % 2;  // Phase3: 翻转
          end
        end

        // pi135: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi135= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi135= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi135= (i + 135) % 2;  // Phase3: 翻转
          end
        end

        // pi136: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi136= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi136= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi136= (i + 136) % 2;  // Phase3: 翻转
          end
        end

        // pi137: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi137= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi137= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi137= (i + 137) % 2;  // Phase3: 翻转
          end
        end

        // pi138: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi138= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi138= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi138= (i + 138) % 2;  // Phase3: 翻转
          end
        end

        // pi139: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi139= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi139= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi139= (i + 139) % 2;  // Phase3: 翻转
          end
        end

        // pi140: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi140= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi140= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi140= (i + 140) % 2;  // Phase3: 翻转
          end
        end

        // pi141: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi141= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi141= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi141= (i + 141) % 2;  // Phase3: 翻转
          end
        end

        // pi142: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi142= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi142= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi142= (i + 142) % 2;  // Phase3: 翻转
          end
        end

        // pi143: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi143= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi143= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi143= (i + 143) % 2;  // Phase3: 翻转
          end
        end

        // pi144: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi144= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi144= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi144= (i + 144) % 2;  // Phase3: 翻转
          end
        end

        // pi145: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi145= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi145= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi145= (i + 145) % 2;  // Phase3: 翻转
          end
        end

        // pi146: 1-bit 三阶段 (稀疏更新)
        if ((i % 4) == 0) begin
          if (i < 170) begin
            pi146= 1'b0;  // Phase1: 全0 (检测SA1)
          end else if (i < 340) begin
            pi146= 1'b1;  // Phase2: 全1 (检测SA0)
          end else begin
            pi146= (i + 146) % 2;  // Phase3: 翻转
          end
        end

      #10;

      if ((i % PRINT_EVERY) == 0) begin
        $display("o_sum=%06x", {po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141});
      end
    end

    $display("o_sum=%06x [final]", {po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141});
    $finish;
  end

  // VCD output
  reg [510:0] dumpfile_name;
  initial begin
    if (!$value$plusargs("DUMPFILE=%s", dumpfile_name)) begin
      $display("Error: No +DUMPFILE argument");
      $finish;
    end
    $display("Dumping VCD to: %s", dumpfile_name);
    $dumpfile(dumpfile_name);
    $dumpvars(0, tb);
  end

  initial begin
    #1;
    $display("FAULT_INJECTED: check_if_force_took_effect");
  end

endmodule
