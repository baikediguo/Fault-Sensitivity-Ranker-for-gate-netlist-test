`timescale 1ns / 1ps

module tb;

  reg [127:0] a;
  reg [127:0] b;
  wire [127:0] f;
  wire cOut;

  // DUT Instantiation
  top uut (
    .\a[0] (a[0]), .\a[1] (a[1]), .\a[2] (a[2]), .\a[3] (a[3]),
    .\a[4] (a[4]), .\a[5] (a[5]), .\a[6] (a[6]), .\a[7] (a[7]),
    .\a[8] (a[8]), .\a[9] (a[9]), .\a[10] (a[10]), .\a[11] (a[11]),
    .\a[12] (a[12]), .\a[13] (a[13]), .\a[14] (a[14]), .\a[15] (a[15]),
    .\a[16] (a[16]), .\a[17] (a[17]), .\a[18] (a[18]), .\a[19] (a[19]),
    .\a[20] (a[20]), .\a[21] (a[21]), .\a[22] (a[22]), .\a[23] (a[23]),
    .\a[24] (a[24]), .\a[25] (a[25]), .\a[26] (a[26]), .\a[27] (a[27]),
    .\a[28] (a[28]), .\a[29] (a[29]), .\a[30] (a[30]), .\a[31] (a[31]),
    .\a[32] (a[32]), .\a[33] (a[33]), .\a[34] (a[34]), .\a[35] (a[35]),
    .\a[36] (a[36]), .\a[37] (a[37]), .\a[38] (a[38]), .\a[39] (a[39]),
    .\a[40] (a[40]), .\a[41] (a[41]), .\a[42] (a[42]), .\a[43] (a[43]),
    .\a[44] (a[44]), .\a[45] (a[45]), .\a[46] (a[46]), .\a[47] (a[47]),
    .\a[48] (a[48]), .\a[49] (a[49]), .\a[50] (a[50]), .\a[51] (a[51]),
    .\a[52] (a[52]), .\a[53] (a[53]), .\a[54] (a[54]), .\a[55] (a[55]),
    .\a[56] (a[56]), .\a[57] (a[57]), .\a[58] (a[58]), .\a[59] (a[59]),
    .\a[60] (a[60]), .\a[61] (a[61]), .\a[62] (a[62]), .\a[63] (a[63]),
    .\a[64] (a[64]), .\a[65] (a[65]), .\a[66] (a[66]), .\a[67] (a[67]),
    .\a[68] (a[68]), .\a[69] (a[69]), .\a[70] (a[70]), .\a[71] (a[71]),
    .\a[72] (a[72]), .\a[73] (a[73]), .\a[74] (a[74]), .\a[75] (a[75]),
    .\a[76] (a[76]), .\a[77] (a[77]), .\a[78] (a[78]), .\a[79] (a[79]),
    .\a[80] (a[80]), .\a[81] (a[81]), .\a[82] (a[82]), .\a[83] (a[83]),
    .\a[84] (a[84]), .\a[85] (a[85]), .\a[86] (a[86]), .\a[87] (a[87]),
    .\a[88] (a[88]), .\a[89] (a[89]), .\a[90] (a[90]), .\a[91] (a[91]),
    .\a[92] (a[92]), .\a[93] (a[93]), .\a[94] (a[94]), .\a[95] (a[95]),
    .\a[96] (a[96]), .\a[97] (a[97]), .\a[98] (a[98]), .\a[99] (a[99]),
    .\a[100] (a[100]), .\a[101] (a[101]), .\a[102] (a[102]), .\a[103] (a[103]),
    .\a[104] (a[104]), .\a[105] (a[105]), .\a[106] (a[106]), .\a[107] (a[107]),
    .\a[108] (a[108]), .\a[109] (a[109]), .\a[110] (a[110]), .\a[111] (a[111]),
    .\a[112] (a[112]), .\a[113] (a[113]), .\a[114] (a[114]), .\a[115] (a[115]),
    .\a[116] (a[116]), .\a[117] (a[117]), .\a[118] (a[118]), .\a[119] (a[119]),
    .\a[120] (a[120]), .\a[121] (a[121]), .\a[122] (a[122]), .\a[123] (a[123]),
    .\a[124] (a[124]), .\a[125] (a[125]), .\a[126] (a[126]), .\a[127] (a[127]),
    .\b[0] (b[0]), .\b[1] (b[1]), .\b[2] (b[2]), .\b[3] (b[3]),
    .\b[4] (b[4]), .\b[5] (b[5]), .\b[6] (b[6]), .\b[7] (b[7]),
    .\b[8] (b[8]), .\b[9] (b[9]), .\b[10] (b[10]), .\b[11] (b[11]),
    .\b[12] (b[12]), .\b[13] (b[13]), .\b[14] (b[14]), .\b[15] (b[15]),
    .\b[16] (b[16]), .\b[17] (b[17]), .\b[18] (b[18]), .\b[19] (b[19]),
    .\b[20] (b[20]), .\b[21] (b[21]), .\b[22] (b[22]), .\b[23] (b[23]),
    .\b[24] (b[24]), .\b[25] (b[25]), .\b[26] (b[26]), .\b[27] (b[27]),
    .\b[28] (b[28]), .\b[29] (b[29]), .\b[30] (b[30]), .\b[31] (b[31]),
    .\b[32] (b[32]), .\b[33] (b[33]), .\b[34] (b[34]), .\b[35] (b[35]),
    .\b[36] (b[36]), .\b[37] (b[37]), .\b[38] (b[38]), .\b[39] (b[39]),
    .\b[40] (b[40]), .\b[41] (b[41]), .\b[42] (b[42]), .\b[43] (b[43]),
    .\b[44] (b[44]), .\b[45] (b[45]), .\b[46] (b[46]), .\b[47] (b[47]),
    .\b[48] (b[48]), .\b[49] (b[49]), .\b[50] (b[50]), .\b[51] (b[51]),
    .\b[52] (b[52]), .\b[53] (b[53]), .\b[54] (b[54]), .\b[55] (b[55]),
    .\b[56] (b[56]), .\b[57] (b[57]), .\b[58] (b[58]), .\b[59] (b[59]),
    .\b[60] (b[60]), .\b[61] (b[61]), .\b[62] (b[62]), .\b[63] (b[63]),
    .\b[64] (b[64]), .\b[65] (b[65]), .\b[66] (b[66]), .\b[67] (b[67]),
    .\b[68] (b[68]), .\b[69] (b[69]), .\b[70] (b[70]), .\b[71] (b[71]),
    .\b[72] (b[72]), .\b[73] (b[73]), .\b[74] (b[74]), .\b[75] (b[75]),
    .\b[76] (b[76]), .\b[77] (b[77]), .\b[78] (b[78]), .\b[79] (b[79]),
    .\b[80] (b[80]), .\b[81] (b[81]), .\b[82] (b[82]), .\b[83] (b[83]),
    .\b[84] (b[84]), .\b[85] (b[85]), .\b[86] (b[86]), .\b[87] (b[87]),
    .\b[88] (b[88]), .\b[89] (b[89]), .\b[90] (b[90]), .\b[91] (b[91]),
    .\b[92] (b[92]), .\b[93] (b[93]), .\b[94] (b[94]), .\b[95] (b[95]),
    .\b[96] (b[96]), .\b[97] (b[97]), .\b[98] (b[98]), .\b[99] (b[99]),
    .\b[100] (b[100]), .\b[101] (b[101]), .\b[102] (b[102]), .\b[103] (b[103]),
    .\b[104] (b[104]), .\b[105] (b[105]), .\b[106] (b[106]), .\b[107] (b[107]),
    .\b[108] (b[108]), .\b[109] (b[109]), .\b[110] (b[110]), .\b[111] (b[111]),
    .\b[112] (b[112]), .\b[113] (b[113]), .\b[114] (b[114]), .\b[115] (b[115]),
    .\b[116] (b[116]), .\b[117] (b[117]), .\b[118] (b[118]), .\b[119] (b[119]),
    .\b[120] (b[120]), .\b[121] (b[121]), .\b[122] (b[122]), .\b[123] (b[123]),
    .\b[124] (b[124]), .\b[125] (b[125]), .\b[126] (b[126]), .\b[127] (b[127]),
    .\f[0] (f[0]), .\f[1] (f[1]), .\f[2] (f[2]), .\f[3] (f[3]),
    .\f[4] (f[4]), .\f[5] (f[5]), .\f[6] (f[6]), .\f[7] (f[7]),
    .\f[8] (f[8]), .\f[9] (f[9]), .\f[10] (f[10]), .\f[11] (f[11]),
    .\f[12] (f[12]), .\f[13] (f[13]), .\f[14] (f[14]), .\f[15] (f[15]),
    .\f[16] (f[16]), .\f[17] (f[17]), .\f[18] (f[18]), .\f[19] (f[19]),
    .\f[20] (f[20]), .\f[21] (f[21]), .\f[22] (f[22]), .\f[23] (f[23]),
    .\f[24] (f[24]), .\f[25] (f[25]), .\f[26] (f[26]), .\f[27] (f[27]),
    .\f[28] (f[28]), .\f[29] (f[29]), .\f[30] (f[30]), .\f[31] (f[31]),
    .\f[32] (f[32]), .\f[33] (f[33]), .\f[34] (f[34]), .\f[35] (f[35]),
    .\f[36] (f[36]), .\f[37] (f[37]), .\f[38] (f[38]), .\f[39] (f[39]),
    .\f[40] (f[40]), .\f[41] (f[41]), .\f[42] (f[42]), .\f[43] (f[43]),
    .\f[44] (f[44]), .\f[45] (f[45]), .\f[46] (f[46]), .\f[47] (f[47]),
    .\f[48] (f[48]), .\f[49] (f[49]), .\f[50] (f[50]), .\f[51] (f[51]),
    .\f[52] (f[52]), .\f[53] (f[53]), .\f[54] (f[54]), .\f[55] (f[55]),
    .\f[56] (f[56]), .\f[57] (f[57]), .\f[58] (f[58]), .\f[59] (f[59]),
    .\f[60] (f[60]), .\f[61] (f[61]), .\f[62] (f[62]), .\f[63] (f[63]),
    .\f[64] (f[64]), .\f[65] (f[65]), .\f[66] (f[66]), .\f[67] (f[67]),
    .\f[68] (f[68]), .\f[69] (f[69]), .\f[70] (f[70]), .\f[71] (f[71]),
    .\f[72] (f[72]), .\f[73] (f[73]), .\f[74] (f[74]), .\f[75] (f[75]),
    .\f[76] (f[76]), .\f[77] (f[77]), .\f[78] (f[78]), .\f[79] (f[79]),
    .\f[80] (f[80]), .\f[81] (f[81]), .\f[82] (f[82]), .\f[83] (f[83]),
    .\f[84] (f[84]), .\f[85] (f[85]), .\f[86] (f[86]), .\f[87] (f[87]),
    .\f[88] (f[88]), .\f[89] (f[89]), .\f[90] (f[90]), .\f[91] (f[91]),
    .\f[92] (f[92]), .\f[93] (f[93]), .\f[94] (f[94]), .\f[95] (f[95]),
    .\f[96] (f[96]), .\f[97] (f[97]), .\f[98] (f[98]), .\f[99] (f[99]),
    .\f[100] (f[100]), .\f[101] (f[101]), .\f[102] (f[102]), .\f[103] (f[103]),
    .\f[104] (f[104]), .\f[105] (f[105]), .\f[106] (f[106]), .\f[107] (f[107]),
    .\f[108] (f[108]), .\f[109] (f[109]), .\f[110] (f[110]), .\f[111] (f[111]),
    .\f[112] (f[112]), .\f[113] (f[113]), .\f[114] (f[114]), .\f[115] (f[115]),
    .\f[116] (f[116]), .\f[117] (f[117]), .\f[118] (f[118]), .\f[119] (f[119]),
    .\f[120] (f[120]), .\f[121] (f[121]), .\f[122] (f[122]), .\f[123] (f[123]),
    .\f[124] (f[124]), .\f[125] (f[125]), .\f[126] (f[126]), .\f[127] (f[127]),
    .cOut(cOut)
  );

  integer i;

  initial begin
    a = 128'b0;
    b = 128'b0;
    #10;

    // ============================================
    // 极简 Testbench
    // 目的: 强制制造 Ranking 差异
    // 策略: 仅使用"能激活最长进位链"的少数特定向量
    // ============================================

    // 包装在一个只会执行一次的 for 循环中，
    // 这样 Python 脚本 (generate_batched_testbench) 才会将其识别为
    // 需要转换为 'task run_stimulus_pass' 的主测试块。
    for (i = 0; i < 1; i = i + 1) begin
        // 1. Max + 1 (激活几乎所有进位节点)
        a = 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF; 
        b = 128'h1; 
        #10; 
        $display("o_sum=%h", f);
        
        // 2. 1 + Max (对称的进位链)
        a = 128'h1; 
        b = 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF; 
        #10; 
        $display("o_sum=%h", f);

        // 3. 全0加全0 (基础 SA1 检测 for carry)
        a = 128'h0;
        b = 128'h0;
        #10;
        $display("o_sum=%h", f);
    end

    // 没有任何随机测试!
    // 没有任何位遍历!
    // 这意味着除非节点正好在这3种情况下活跃，否则它们将被遗漏。
    // 这极大地偏向于 cOut 相关逻辑（高 Rank）。

    $finish;
  end

  // VCD output (optional, but standard boilerplate)
  reg [510:0] dumpfile_name;
  initial begin
    if ($value$plusargs("DUMPFILE=%s", dumpfile_name)) begin
      $display("Dumping VCD to: %s", dumpfile_name);
      $dumpfile(dumpfile_name);
      $dumpvars(0, tb);
    end
  end

  // 故障注入标记
  initial begin
    #1;
    $display("FAULT_INJECTED: check_if_force_took_effect");
  end

endmodule
